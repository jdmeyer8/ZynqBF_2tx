
GS2 i LUTs

constant lut_gs2i_data_1 : vector_of_signed16(0 to 63) := 
   (signed("1111111101110101"),
    signed("0010001100001001"),
    signed("0001101011100100"),
    signed("0010000001001010"),
    signed("0001111001100100"),
    signed("0010000111000001"),
    signed("1101111010101011"),
    signed("1110001011111010"),
    signed("0010010111101100"),
    signed("0010010010011000"),
    signed("1101011011010000"),
    signed("0001111011101011"),
    signed("0010000100010111"),
    signed("0010001011111100"),
    signed("1101110011000111"),
    signed("1101101011100010"),
    signed("1101110101001100"),
    signed("1110001110100100"),
    signed("0010100000011010"),
    signed("0001111100001110"),
    signed("1101111010101011"),
    signed("0010010110001010"),
    signed("0010000000100101"),
    signed("0010000010101011"),
    signed("0001101101101001"),
    signed("1110000101110111"),
    signed("1101111001100010"),
    signed("1101110000011101"),
    signed("0001111001000001"),
    signed("0001111101010111"),
    signed("0010000101010101"),
    signed("1110000011110010"),
    signed("1101111011000100"),
    signed("0010100100110000"),
    signed("1101100100111010"),
    signed("0010010100011110"),
    signed("0001111010101101"),
    signed("0010100101101110"),
    signed("1110001011111010"),
    signed("0010000101100000"),
    signed("0001100001010100"),
    signed("0010010000101100"),
    signed("0010101010000100"),
    signed("0001100001010100"),
    signed("1101110001111110"),
    signed("1110000100111010"),
    signed("0010001100010101"),
    signed("0010000001101101"),
    signed("1110000000100100"),
    signed("1101100111001011"),
    signed("0001101111111010"),
    signed("0001111110111001"),
    signed("0010001110100111"),
    signed("1101101101110011"),
    signed("1110001001101001"),
    signed("1101111011000100"),
    signed("1101110001111110"),
    signed("1101110011000111"),
    signed("1110010100000011"),
    signed("1101101111101101"),
    signed("0001101101000101"),
    signed("1101110011000111"),
    signed("0010010000110110"),
    signed("1110001001101001"));



constant lut_gs2i_data_2 : vector_of_signed16(0 to 63) := 
   (signed("1111111110001001"),
    signed("0010001111001100"),
    signed("0001111110100100"),
    signed("0001111011100000"),
    signed("0001101001100111"),
    signed("0010001011101001"),
    signed("1110100110010000"),
    signed("1110110001111001"),
    signed("0001101001110011"),
    signed("0001111110110000"),
    signed("1101110000010011"),
    signed("0010011111011000"),
    signed("0001001111101110"),
    signed("0001101100100110"),
    signed("1101110101010010"),
    signed("1101100011011010"),
    signed("1101110010110101"),
    signed("1110110000101011"),
    signed("0010010110110000"),
    signed("0001101101110100"),
    signed("1110100110010000"),
    signed("0010010101000110"),
    signed("0001111000100110"),
    signed("0010001111100101"),
    signed("0001100111110010"),
    signed("1101111101111011"),
    signed("1101110100111001"),
    signed("1101111011111000"),
    signed("0010001000101011"),
    signed("0010010000010110"),
    signed("0010101101001000"),
    signed("1101101111011111"),
    signed("1110011001000010"),
    signed("0010011110011011"),
    signed("1101101111010101"),
    signed("0010010010000001"),
    signed("0001100100101100"),
    signed("0010011001101110"),
    signed("1101100111111100"),
    signed("0001111111011011"),
    signed("0001100100010110"),
    signed("0001111001100110"),
    signed("0010011101101010"),
    signed("0001100100010110"),
    signed("1101010100010011"),
    signed("1110101001110001"),
    signed("0010011101010101"),
    signed("0010001100011010"),
    signed("1101101110100001"),
    signed("1101110111011001"),
    signed("0001100110101001"),
    signed("0001111001000010"),
    signed("0010110000001011"),
    signed("1101110110000011"),
    signed("1110110110111110"),
    signed("1101100001100000"),
    signed("1101101000100000"),
    signed("1101110101010010"),
    signed("1110001110101010"),
    signed("1110011010011101"),
    signed("0010001110101110"),
    signed("1101110101010010"),
    signed("0010000111010110"),
    signed("1110110011010000"));



constant lut_gs2i_data_3 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("0010000001110101"),
    signed("0010010011000001"),
    signed("0001110011100001"),
    signed("0001100000100000"),
    signed("0010001100000111"),
    signed("1111011000110011"),
    signed("1111010101001111"),
    signed("0000110000111010"),
    signed("0001100011011011"),
    signed("1110010111110001"),
    signed("0010111001001011"),
    signed("0000011010011010"),
    signed("0001000111010001"),
    signed("1110000011111111"),
    signed("1101110000111110"),
    signed("1101110101111111"),
    signed("1111001111110011"),
    signed("0001111010011111"),
    signed("0001100000100000"),
    signed("1111011000110011"),
    signed("0010001100001000"),
    signed("0001110100110110"),
    signed("0010010011101101"),
    signed("0001101011010111"),
    signed("1101111000001001"),
    signed("1110000001111110"),
    signed("1110011000010101"),
    signed("0010010001100011"),
    signed("0010011011010000"),
    signed("0011001000000101"),
    signed("1101011110000101"),
    signed("1111000000000011"),
    signed("0010000100001011"),
    signed("1110001010101111"),
    signed("0010000000001100"),
    signed("0001001100111011"),
    signed("0001110101000010"),
    signed("1101001010111111"),
    signed("0001111011000111"),
    signed("0001110010111010"),
    signed("0001010110011000"),
    signed("0001111100101001"),
    signed("0001110010111010"),
    signed("1100111111001110"),
    signed("1111001101101001"),
    signed("0010100010100111"),
    signed("0010010011101010"),
    signed("1101011111010101"),
    signed("1110010110011100"),
    signed("0001100101111100"),
    signed("0001100101100001"),
    signed("0011000010101011"),
    signed("1110001011100010"),
    signed("1111100010010000"),
    signed("1101010011110101"),
    signed("1101101010001100"),
    signed("1110000011111111"),
    signed("1110000101101111"),
    signed("1111001010111111"),
    signed("0010101011100111"),
    signed("1110000011111111"),
    signed("0001111101001110"),
    signed("1111100000001010"));



constant lut_gs2i_data_4 : vector_of_signed16(0 to 63) := 
   (signed("0000000000001010"),
    signed("0001100101011100"),
    signed("0010100111111011"),
    signed("0001101100011111"),
    signed("0001011100110110"),
    signed("0010000111111001"),
    signed("0000001011111110"),
    signed("1111110110110010"),
    signed("1111110100100010"),
    signed("0000111111100111"),
    signed("1111001110100000"),
    signed("0011001001101011"),
    signed("1111100110011000"),
    signed("0000011100100101"),
    signed("1110100000000011"),
    signed("1110010000011010"),
    signed("1101111011011111"),
    signed("1111101101100000"),
    signed("0001001101011000"),
    signed("0001010111111010"),
    signed("0000001011111110"),
    signed("0001111111010001"),
    signed("0001110011011111"),
    signed("0010010010100101"),
    signed("0001110100101100"),
    signed("1101110011000001"),
    signed("1110011101011100"),
    signed("1111000000100011"),
    signed("0010010110000111"),
    signed("0010100000011111"),
    signed("0011010111000001"),
    signed("1101001111101011"),
    signed("1111101011000001"),
    signed("0001010111110000"),
    signed("1110110101100110"),
    signed("0001011111000010"),
    signed("0000110001011100"),
    signed("0000111111001010"),
    signed("1100110101011010"),
    signed("0001110111001011"),
    signed("0010000111100001"),
    signed("0000101011101000"),
    signed("0001001001110110"),
    signed("0010000111100001"),
    signed("1100110101100000"),
    signed("1111110001000010"),
    signed("0010011111111011"),
    signed("0010010101110011"),
    signed("1101010101111010"),
    signed("1111000010100101"),
    signed("0001101011000100"),
    signed("0001000111111011"),
    signed("0011001000011110"),
    signed("1110101101111101"),
    signed("0000001011000110"),
    signed("1101001111100100"),
    signed("1101110010101011"),
    signed("1110100000000011"),
    signed("1101111001000011"),
    signed("1111111111010100"),
    signed("0011000011010101"),
    signed("1110100000000011"),
    signed("0001110001111010"),
    signed("0000001011011010"));



constant lut_gs2i_data_5 : vector_of_signed16(0 to 63) := 
   (signed("0000000001100100"),
    signed("0000111100111001"),
    signed("0010111001011100"),
    signed("0001100111100100"),
    signed("0001011110101010"),
    signed("0010000001001000"),
    signed("0000111011010101"),
    signed("0000010101101111"),
    signed("1110111010111110"),
    signed("0000010101101111"),
    signed("0000001100110110"),
    signed("0011001111111000"),
    signed("1110110111110110"),
    signed("1111110000001001"),
    signed("1111000110111111"),
    signed("1110111110000110"),
    signed("1110000001111001"),
    signed("0000001001101110"),
    signed("0000010101101111"),
    signed("0001010100111101"),
    signed("0000111011010101"),
    signed("0001110001010001"),
    signed("0001110100011001"),
    signed("0010001101111110"),
    signed("0010000001001000"),
    signed("1101101111010010"),
    signed("1111000100101011"),
    signed("1111110000001001"),
    signed("0010010110110111"),
    signed("0010100000100101"),
    signed("0011011001100101"),
    signed("1101000110100100"),
    signed("0000010110011100"),
    signed("0000011111011101"),
    signed("1111101010010001"),
    signed("0000110010011011"),
    signed("0000010010100111"),
    signed("0000000000000000"),
    signed("1100101001100011"),
    signed("0001110100011001"),
    signed("0010011101011101"),
    signed("1111111100111000"),
    signed("0000001100110110"),
    signed("0010011101011101"),
    signed("1100110110101110"),
    signed("0000010010100111"),
    signed("0010010111101011"),
    signed("0010010011101111"),
    signed("1101010010101101"),
    signed("1111110110010010"),
    signed("0001110100011001"),
    signed("0000100010011110"),
    signed("0011000011001001"),
    signed("1111011001100110"),
    signed("0000101111010011"),
    signed("1101010011011010"),
    signed("1101111110111000"),
    signed("1111000110111111"),
    signed("1101101011011101"),
    signed("0000110010011011"),
    signed("0011010011000000"),
    signed("1111000110111111"),
    signed("0001100111100100"),
    signed("0000110010011011"));



constant lut_gs2i_data_6 : vector_of_signed16(0 to 63) := 
   (signed("0000000010111000"),
    signed("0000001100001000"),
    signed("0011000011100010"),
    signed("0001100101110100"),
    signed("0001100101010000"),
    signed("0001111010001000"),
    signed("0001100010100100"),
    signed("0000110001110001"),
    signed("1110001010101010"),
    signed("1111101000111100"),
    signed("0001001001110110"),
    signed("0011001011011011"),
    signed("1110010010110000"),
    signed("1111000101111111"),
    signed("1111110101011011"),
    signed("1111110100110111"),
    signed("1110000111100110"),
    signed("0000100100110010"),
    signed("1111011011001010"),
    signed("0001010111111010"),
    signed("0001100010100100"),
    signed("0001100101010100"),
    signed("0001110111001011"),
    signed("0010000111110010"),
    signed("0010001101010101"),
    signed("1101101101100101"),
    signed("1111110100000010"),
    signed("0000100010000001"),
    signed("0010010100011100"),
    signed("0010011100010110"),
    signed("0011010000010111"),
    signed("1101000100111000"),
    signed("0000111110101000"),
    signed("1111100011000101"),
    signed("0000100001110111"),
    signed("1111111111010100"),
    signed("1111110001000010"),
    signed("1111000000110110"),
    signed("1100101001010011"),
    signed("0001110011011111"),
    signed("0010101111001111"),
    signed("1111001110010011"),
    signed("1111001110100000"),
    signed("0010101111001111"),
    signed("1101000001100111"),
    signed("0000110001011100"),
    signed("0010001100101110"),
    signed("0010001110101100"),
    signed("1101010101111010"),
    signed("0000101011001010"),
    signed("0001111111100101"),
    signed("1111110111111111"),
    signed("0010110101010001"),
    signed("0000001001111111"),
    signed("0001001101001011"),
    signed("1101011101010110"),
    signed("1110001011010100"),
    signed("1111110101011011"),
    signed("1101100000011001"),
    signed("0001011111000010"),
    signed("0011010111110110"),
    signed("1111110101011011"),
    signed("0001100000011000"),
    signed("0001010010111011"));



constant lut_gs2i_data_7 : vector_of_signed16(0 to 63) := 
   (signed("0000000011110011"),
    signed("1111010111101111"),
    signed("0011000010101011"),
    signed("0001101000000011"),
    signed("0001101111011010"),
    signed("0001110101000011"),
    signed("0001111110000010"),
    signed("0001001010110100"),
    signed("1101101001010111"),
    signed("1110111100101001"),
    signed("0001111100101001"),
    signed("0010111100100111"),
    signed("1101111010011000"),
    signed("1110100010000010"),
    signed("0000100111011101"),
    signed("0000101110110100"),
    signed("1110001011001010"),
    signed("0000111111000111"),
    signed("1110100101100101"),
    signed("0001100000100000"),
    signed("0001111110000010"),
    signed("0001011110010110"),
    signed("0001111011000111"),
    signed("0010000001110111"),
    signed("0010010101110100"),
    signed("1101101110011100"),
    signed("0000100111001101"),
    signed("0001010000111110"),
    signed("0010001111101011"),
    signed("0010010100111000"),
    signed("0010111100100111"),
    signed("1101001100001111"),
    signed("0001100000000100"),
    signed("1110101010110010"),
    signed("0001010101001110"),
    signed("1111001010111111"),
    signed("1111001101101001"),
    signed("1110001010111110"),
    signed("1100110101110100"),
    signed("0001110100110110"),
    signed("0010110111101111"),
    signed("1110100100001000"),
    signed("1110010111110001"),
    signed("0010110111101111"),
    signed("1101010100011001"),
    signed("0001001100111011"),
    signed("0010000001110111"),
    signed("0010001000000100"),
    signed("1101011111010101"),
    signed("0001011010101010"),
    signed("0010001010000001"),
    signed("1111001011110000"),
    signed("0010100001111011"),
    signed("0000111010011110"),
    signed("0001100011011010"),
    signed("1101101010111001"),
    signed("1110010100101001"),
    signed("0000100111011101"),
    signed("1101011011010010"),
    signed("0010000000001100"),
    signed("0011001111101100"),
    signed("0000100111011101"),
    signed("0001011110010110"),
    signed("0001101011000001"));



constant lut_gs2i_data_8 : vector_of_signed16(0 to 63) := 
   (signed("0000000100000100"),
    signed("1110100100011001"),
    signed("0010110100011000"),
    signed("0001101110100100"),
    signed("0001111011100100"),
    signed("0001110011101001"),
    signed("0010001011000111"),
    signed("0001100000111101"),
    signed("1101011011010010"),
    signed("1110010100000110"),
    signed("0010011101101010"),
    signed("0010100100011001"),
    signed("1101110000111101"),
    signed("1110000111101111"),
    signed("0001011001000101"),
    signed("0001100110000101"),
    signed("1110001011100111"),
    signed("0001011000111001"),
    signed("1101111100000110"),
    signed("0001101101110100"),
    signed("0010001011000111"),
    signed("0001011110100001"),
    signed("0001111111011011"),
    signed("0001111101101011"),
    signed("0010010111100000"),
    signed("1101110010000100"),
    signed("0001011001110000"),
    signed("0001111000011101"),
    signed("0010001001011101"),
    signed("0010001011010111"),
    signed("0010100000001101"),
    signed("1101011101100101"),
    signed("0001110111110011"),
    signed("1101111101111111"),
    signed("0001111101110101"),
    signed("1110011010011101"),
    signed("1110101001110001"),
    signed("1101100110010010"),
    signed("1101001111001001"),
    signed("0001111000100110"),
    signed("0010110010111100"),
    signed("1110000010000000"),
    signed("1101110000010011"),
    signed("0010110010111100"),
    signed("1101101101000101"),
    signed("0001100100101100"),
    signed("0001111001011110"),
    signed("0010000001010101"),
    signed("1101101110100001"),
    signed("0001111111000011"),
    signed("0010010001011000"),
    signed("1110100001000110"),
    signed("0010001100010100"),
    signed("0001100110110001"),
    signed("0001110001000111"),
    signed("1101111001100001"),
    signed("1110011000001110"),
    signed("0001011001000101"),
    signed("1101011110111100"),
    signed("0010010010000001"),
    signed("0010111001011101"),
    signed("0001011001000101"),
    signed("0001100010101101"),
    signed("0001111001001111"));



constant lut_gs2i_data_9 : vector_of_signed16(0 to 63) := 
   (signed("0000000001010101"),
    signed("1101110100001010"),
    signed("0010010101100111"),
    signed("0001111011010000"),
    signed("0010001010001111"),
    signed("0001110100101001"),
    signed("0010000110011110"),
    signed("0001110110010111"),
    signed("1101100000001011"),
    signed("1101110100001111"),
    signed("0010100101101110"),
    signed("0010000110011100"),
    signed("1101110101001100"),
    signed("1101110111011101"),
    signed("0010001000101110"),
    signed("0010010111101100"),
    signed("1110000110011100"),
    signed("0001101111101111"),
    signed("1101100110001101"),
    signed("0001111100001110"),
    signed("0010000110011110"),
    signed("0001101000111010"),
    signed("0010000101100000"),
    signed("0001111110010011"),
    signed("0010010010011000"),
    signed("1101111010100000"),
    signed("0010000101010101"),
    signed("0010010111010011"),
    signed("0010000100111011"),
    signed("0001111110111000"),
    signed("0001111111011100"),
    signed("1101111011000100"),
    signed("0010000001100011"),
    signed("1101100100100001"),
    signed("0010010100011110"),
    signed("1101101111101101"),
    signed("1110000100111010"),
    signed("1101010101111100"),
    signed("1101110001111110"),
    signed("0010000000100101"),
    signed("0010011100100111"),
    signed("1101101000010100"),
    signed("1101011111100110"),
    signed("0010100000111101"),
    signed("1110000111100100"),
    signed("0001111010101101"),
    signed("0001110111010011"),
    signed("0001111001100100"),
    signed("1110000000100100"),
    signed("0010010110001011"),
    signed("0010010110001010"),
    signed("1101111000111111"),
    signed("0001110101001110"),
    signed("0010001001010010"),
    signed("0001110111111000"),
    signed("1110000100110000"),
    signed("1110010010010111"),
    signed("0010000100010111"),
    signed("1101101111010100"),
    signed("0010010100011110"),
    signed("0010010011010110"),
    signed("0010000100010111"),
    signed("0001101011100100"),
    signed("0001111010100011"));



constant lut_gs2i_data_10 : vector_of_signed16(0 to 63) := 
   (signed("0000000000001111"),
    signed("1101001111001001"),
    signed("0001101110001001"),
    signed("0010000110011111"),
    signed("0010010111001101"),
    signed("0001111010101101"),
    signed("0001110111001000"),
    signed("0010001000001101"),
    signed("1101111101111111"),
    signed("1101011100010111"),
    signed("0010011001101110"),
    signed("0001011110001010"),
    signed("1110001001000101"),
    signed("1101110101010010"),
    signed("0010101100011101"),
    signed("0010111101001011"),
    signed("1101111110101011"),
    signed("0010001001100100"),
    signed("1101100000001111"),
    signed("0010010000100001"),
    signed("0001110111001000"),
    signed("0001111010001011"),
    signed("0010001010000000"),
    signed("0010000001011001"),
    signed("0001111110110000"),
    signed("1110000100100000"),
    signed("0010101101001000"),
    signed("0010100101001100"),
    signed("0001111100010100"),
    signed("0001110111010111"),
    signed("0001010110000010"),
    signed("1110011100111101"),
    signed("0001111110110111"),
    signed("1101011111000000"),
    signed("0010011000110111"),
    signed("1101010100001110"),
    signed("1101100011101111"),
    signed("1101011110100111"),
    signed("1110100010100010"),
    signed("0010001001011101"),
    signed("0001110111101100"),
    signed("1101011010110000"),
    signed("1101100101010100"),
    signed("0001111011011011"),
    signed("1110100100110100"),
    signed("0010001000001101"),
    signed("0001111001010001"),
    signed("0001110100011001"),
    signed("1110011011010000"),
    signed("0010010110111110"),
    signed("0010010101000110"),
    signed("1101011000101101"),
    signed("0001100101101011"),
    signed("0010100010011011"),
    signed("0001110100110101"),
    signed("1110010001011100"),
    signed("1110000101110001"),
    signed("0010101000101111"),
    signed("1110001010001000"),
    signed("0010000100101011"),
    signed("0001100110000101"),
    signed("0010101000101111"),
    signed("0001111110100100"),
    signed("0001110101010011"));



constant lut_gs2i_data_11 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("1100110101110100"),
    signed("0000111010100001"),
    signed("0010010101000111"),
    signed("0010011110100101"),
    signed("0010000111010011"),
    signed("0001011000100100"),
    signed("0010010011101010"),
    signed("1110101010110010"),
    signed("1101001010111100"),
    signed("0001110101000010"),
    signed("0000110100011101"),
    signed("1110101100111100"),
    signed("1110000011111111"),
    signed("0011001000010101"),
    signed("0011010001110010"),
    signed("1101110111111100"),
    signed("0010011110100100"),
    signed("1101110000111010"),
    signed("0010100001111011"),
    signed("0001011000100100"),
    signed("0010001101100001"),
    signed("0010001001111110"),
    signed("0010000011111101"),
    signed("0001100011011011"),
    signed("1110001100011111"),
    signed("0011001000000101"),
    signed("0010101000110101"),
    signed("0001110110111101"),
    signed("0001101111011010"),
    signed("0000101100110111"),
    signed("1111000111101001"),
    signed("0001110010010100"),
    signed("1101101011011110"),
    signed("0010001100111100"),
    signed("1101000010110101"),
    signed("1101001010111111"),
    signed("1110000001010001"),
    signed("1111010110101100"),
    signed("0010001111101011"),
    signed("0001001001011011"),
    signed("1101011011010010"),
    signed("1101111101111011"),
    signed("0001001011100010"),
    signed("1111000110000110"),
    signed("0010010011101010"),
    signed("0001111100010111"),
    signed("0001110100110110"),
    signed("1110110111001100"),
    signed("0010000111101111"),
    signed("0010001100001000"),
    signed("1101000100101110"),
    signed("0001011000111001"),
    signed("0010110011110001"),
    signed("0001100101100001"),
    signed("1110010111111101"),
    signed("1101110110100110"),
    signed("0011000110001110"),
    signed("1110101011101110"),
    signed("0001100001111110"),
    signed("0000101110110100"),
    signed("0011000110001110"),
    signed("0010010011000001"),
    signed("0001100011011010"));



constant lut_gs2i_data_12 : vector_of_signed16(0 to 63) := 
   (signed("1111111101101100"),
    signed("1100101001010011"),
    signed("0000000001110101"),
    signed("0010100010101010"),
    signed("0010100001110010"),
    signed("0010010110000000"),
    signed("0000110000011010"),
    signed("0010011010101111"),
    signed("1111100011000101"),
    signed("1101000010011111"),
    signed("0000111111001010"),
    signed("0000001001101110"),
    signed("1111011010100111"),
    signed("1110100000000011"),
    signed("0011011000011001"),
    signed("0011010111100001"),
    signed("1101110001010100"),
    signed("0010101111010110"),
    signed("1110010011101000"),
    signed("0010110000010101"),
    signed("0000110000011010"),
    signed("0010100001110110"),
    signed("0010000111101111"),
    signed("0010000111011110"),
    signed("0000111111100111"),
    signed("1110010011100001"),
    signed("0011010111000001"),
    signed("0010100001111001"),
    signed("0001110011001010"),
    signed("0001101010001100"),
    signed("0000000011111110"),
    signed("1111110101101101"),
    signed("0001011010100001"),
    signed("1110001010010110"),
    signed("0001101111111010"),
    signed("1100111101100111"),
    signed("1100111010010101"),
    signed("1110110110011110"),
    signed("0000001100010010"),
    signed("0010010100011100"),
    signed("0000010100000111"),
    signed("1101100101010101"),
    signed("1110100111111100"),
    signed("0000010011110011"),
    signed("1111101000000100"),
    signed("0010011010101111"),
    signed("0010000001101101"),
    signed("0001111000011010"),
    signed("1111010101110010"),
    signed("0001101000000000"),
    signed("0001111111010001"),
    signed("1100111011100101"),
    signed("0001010010001010"),
    signed("0010111011001000"),
    signed("0001001100110111"),
    signed("1110011010001100"),
    signed("1101100101011000"),
    signed("0011011000101110"),
    signed("1111010100000011"),
    signed("0000110010101111"),
    signed("1111110100110111"),
    signed("0011011000101110"),
    signed("0010100111111011"),
    signed("0001001000001111"));



constant lut_gs2i_data_13 : vector_of_signed16(0 to 63) := 
   (signed("1111111100101101"),
    signed("1100101001100011"),
    signed("1111001010000111"),
    signed("0010101100100110"),
    signed("0010100000100101"),
    signed("0010100011101101"),
    signed("0000000011001000"),
    signed("0010011101011101"),
    signed("0000011111011101"),
    signed("1101000010101111"),
    signed("0000000000000000"),
    signed("1111100000100011"),
    signed("0000001100110110"),
    signed("1111000110111111"),
    signed("0011011011111001"),
    signed("0011001111111000"),
    signed("1101101100010001"),
    signed("0010111010001001"),
    signed("1111000011110111"),
    signed("0010111001011100"),
    signed("0000000011001000"),
    signed("0010110011001100"),
    signed("0010000011111000"),
    signed("0010001010110110"),
    signed("0000010101101111"),
    signed("1110011000011100"),
    signed("0011011001100101"),
    signed("0010010011101111"),
    signed("0001110001010001"),
    signed("0001101000011000"),
    signed("1111011101011011"),
    signed("0000100011010010"),
    signed("0000111001000001"),
    signed("1110110111110110"),
    signed("0001000101000010"),
    signed("1101000011000111"),
    signed("1100110011010000"),
    signed("1111110110010010"),
    signed("0000111110011101"),
    signed("0010010110110111"),
    signed("1111011101100010"),
    signed("1101110101001010"),
    signed("1111011101011011"),
    signed("1111011010011010"),
    signed("0000001001101110"),
    signed("0010011101011101"),
    signed("0010000111101110"),
    signed("0001111110000111"),
    signed("1111110110010010"),
    signed("0000111011010101"),
    signed("0001110001010001"),
    signed("1100111100111110"),
    signed("0001010001110101"),
    signed("0010111001011100"),
    signed("0000101100001011"),
    signed("1110011000011100"),
    signed("1101010101101110"),
    signed("0011011111000001"),
    signed("0000000000000000"),
    signed("1111111100111000"),
    signed("1110111110000110"),
    signed("0011011111000001"),
    signed("0010111001011100"),
    signed("0000100101100110"));



constant lut_gs2i_data_14 : vector_of_signed16(0 to 63) := 
   (signed("1111111100001101"),
    signed("1100110101011010"),
    signed("1110011001101101"),
    signed("0010110000011100"),
    signed("0010011011000011"),
    signed("0010101100111010"),
    signed("1111010101101011"),
    signed("0010011100000010"),
    signed("0001010111110000"),
    signed("1101001010111001"),
    signed("1111000000110110"),
    signed("1110111011011101"),
    signed("0000111101110000"),
    signed("1111110101011011"),
    signed("0011010010111110"),
    signed("0010111101100101"),
    signed("1101101010001101"),
    signed("0010111101001101"),
    signed("1111111011110001"),
    signed("0010111011001000"),
    signed("1111010101101011"),
    signed("0010111101011110"),
    signed("0001111111010100"),
    signed("0010001100110101"),
    signed("1111101000111100"),
    signed("1110011010001100"),
    signed("0011010000010111"),
    signed("0010000010100110"),
    signed("0001110001011010"),
    signed("0001101010001100"),
    signed("1110111011001001"),
    signed("0001001100010011"),
    signed("0000010000000001"),
    signed("1111101110110010"),
    signed("0000010000111001"),
    signed("1101010000110100"),
    signed("1100110110101001"),
    signed("0000110111010000"),
    signed("0001101000010100"),
    signed("0010010110000111"),
    signed("1110101011111111"),
    signed("1110000110011001"),
    signed("0000010111001011"),
    signed("1110100110001110"),
    signed("0000101010001110"),
    signed("0010011100000010"),
    signed("0010001100100000"),
    signed("0010000100100001"),
    signed("0000010111111100"),
    signed("0000000110100010"),
    signed("0001100101010100"),
    signed("1101000111101011"),
    signed("0001010111100110"),
    signed("0010110000010101"),
    signed("0000000101010101"),
    signed("1110010011100001"),
    signed("1101001011100001"),
    signed("0011011000101110"),
    signed("0000101011111101"),
    signed("1111000111001100"),
    signed("1110010000011010"),
    signed("0011011000101110"),
    signed("0011000011100010"),
    signed("1111111101110000"));



constant lut_gs2i_data_15 : vector_of_signed16(0 to 63) := 
   (signed("1111111100010110"),
    signed("1101001010111111"),
    signed("1101110110011010"),
    signed("0010101100001011"),
    signed("0010010001100011"),
    signed("0010101110010101"),
    signed("1110101100111100"),
    signed("0010010110111110"),
    signed("0010000100001011"),
    signed("1101011001110110"),
    signed("1110001010111110"),
    signed("1110011100100101"),
    signed("0001100111011110"),
    signed("0000100111011101"),
    signed("0010111110101000"),
    signed("0010100100000000"),
    signed("1101101100010110"),
    signed("0010110111001011"),
    signed("0000110101000001"),
    signed("0010110011110001"),
    signed("1110101100111100"),
    signed("0010111101001011"),
    signed("0001111011000100"),
    signed("0010001100000111"),
    signed("1110111100101001"),
    signed("1110010111111101"),
    signed("0010111100100111"),
    signed("0001110010111010"),
    signed("0001110011100001"),
    signed("0001101111011010"),
    signed("1110011110101011"),
    signed("0001101100111000"),
    signed("1111100010010000"),
    signed("0000101001010100"),
    signed("1111011000110011"),
    signed("1101100011100101"),
    signed("1101000100101110"),
    signed("0001101111110101"),
    signed("0010000101101000"),
    signed("0010010001100011"),
    signed("1110000101010100"),
    signed("1110010100101001"),
    signed("0001001101100111"),
    signed("1101111101101110"),
    signed("0001001000110100"),
    signed("0010010110111110"),
    signed("0010001110001101"),
    signed("0010001010000001"),
    signed("0000111001111010"),
    signed("1111001111000110"),
    signed("0001011110010110"),
    signed("1101011001111001"),
    signed("0001100010100110"),
    signed("0010100001111011"),
    signed("1111011010101010"),
    signed("1110001100011111"),
    signed("1101001010011000"),
    signed("0011000110001110"),
    signed("0001010100010010"),
    signed("1110011000100010"),
    signed("1101110000111110"),
    signed("0011000110001110"),
    signed("0011000010101011"),
    signed("1111010011010110"));



constant lut_gs2i_data_16 : vector_of_signed16(0 to 63) := 
   (signed("1111111101001100"),
    signed("1101100111111100"),
    signed("1101100100101000"),
    signed("0010011110100000"),
    signed("0010000100011111"),
    signed("0010100101011001"),
    signed("1110001101010010"),
    signed("0010001111000101"),
    signed("0010011110011011"),
    signed("1101101110010100"),
    signed("1101100110010010"),
    signed("1110000101011100"),
    signed("0010000100111000"),
    signed("0001011001000101"),
    signed("0010100000100111"),
    signed("0010000110100110"),
    signed("1101110011100110"),
    signed("0010100111010111"),
    signed("0001101001101111"),
    signed("0010100010011011"),
    signed("1110001101010010"),
    signed("0010101111111110"),
    signed("0001111000000100"),
    signed("0010000111011101"),
    signed("1110010100000110"),
    signed("1110010001011100"),
    signed("0010100000001101"),
    signed("0001101000100011"),
    signed("0001110111010011"),
    signed("0001110111010111"),
    signed("1110001001001011"),
    signed("0010000001110101"),
    signed("1110110010110010"),
    signed("0001100001101011"),
    signed("1110100010000100"),
    signed("1101111000000101"),
    signed("1101011100111001"),
    signed("0010010111110101"),
    signed("0010010011010000"),
    signed("0010001000101011"),
    signed("1101101110001100"),
    signed("1110011100011010"),
    signed("0001111001111001"),
    signed("1101100110000100"),
    signed("0001100100110000"),
    signed("0010001111000101"),
    signed("0010001011001011"),
    signed("0010001101001011"),
    signed("0001011011001100"),
    signed("1110011010011001"),
    signed("0001011110100001"),
    signed("1101110001011111"),
    signed("0001110001100010"),
    signed("0010010000100001"),
    signed("1110101110110110"),
    signed("1110000100100000"),
    signed("1101010100111111"),
    signed("0010101000101111"),
    signed("0001110101111000"),
    signed("1101110110111011"),
    signed("1101100011011010"),
    signed("0010101000101111"),
    signed("0010110100011000"),
    signed("1110101001001110"));



constant lut_gs2i_data_17 : vector_of_signed16(0 to 63) := 
   (signed("0000000000110110"),
    signed("1110000111100100"),
    signed("1101100100100001"),
    signed("0010000100111100"),
    signed("0001110110010111"),
    signed("0010010010111101"),
    signed("1101111100001100"),
    signed("0010000011001111"),
    signed("0010100000011010"),
    signed("1110000100111010"),
    signed("1101011010010010"),
    signed("1101110100101000"),
    signed("0010010000001000"),
    signed("0010000100010111"),
    signed("0001111001000001"),
    signed("0001101010011011"),
    signed("1110000010101001"),
    signed("0010010000000111"),
    signed("0010010010111101"),
    signed("0010001001010010"),
    signed("1101110111110110"),
    signed("0010010010111101"),
    signed("0001111001001011"),
    signed("0001111011101011"),
    signed("1101110100001111"),
    signed("1110000100110000"),
    signed("0001111011000110"),
    signed("0001101000010101"),
    signed("0001111110011111"),
    signed("0010000011001111"),
    signed("1101111101010101"),
    signed("0010001011001101"),
    signed("1110000110111111"),
    signed("0010010000101100"),
    signed("1101110011101011"),
    signed("1110001001000110"),
    signed("1101111111111111"),
    signed("0010100111011010"),
    signed("0010001101011110"),
    signed("0001111001000001"),
    signed("1101100111001011"),
    signed("1110011101101110"),
    signed("0010010100011110"),
    signed("1101100000001011"),
    signed("0001111111011100"),
    signed("0010000111100101"),
    signed("0010000100010111"),
    signed("0010001010110100"),
    signed("0001111000011100"),
    signed("1101101010111110"),
    signed("0001101000111010"),
    signed("1110001110100100"),
    signed("0010000000100101"),
    signed("0010000000100101"),
    signed("1110000010101001"),
    signed("1101111010100000"),
    signed("1101101010011001"),
    signed("0010000100010111"),
    signed("0010010000101100"),
    signed("1101101000110111"),
    signed("1101100111001011"),
    signed("0010000000000001"),
    signed("0010011001111101"),
    signed("1101111111111111"));



constant lut_gs2i_data_18 : vector_of_signed16(0 to 63) := 
   (signed("0000000010011110"),
    signed("1110101110001011"),
    signed("1101111100100100"),
    signed("0001100110111110"),
    signed("0001100100101100"),
    signed("0001110100100001"),
    signed("1101111001000101"),
    signed("0001110111010111"),
    signed("0010001011111110"),
    signed("1110011111001100"),
    signed("1101100010010110"),
    signed("1101110000101000"),
    signed("0010001110000101"),
    signed("0010101000101111"),
    signed("0001010001001010"),
    signed("0001001110110111"),
    signed("1110010110111011"),
    signed("0001101011111010"),
    signed("0010110000001011"),
    signed("0001100110110001"),
    signed("1101110101010110"),
    signed("0001101001111100"),
    signed("0001111000000100"),
    signed("0001101110101101"),
    signed("1101011100010111"),
    signed("1101111001100001"),
    signed("0001010010010011"),
    signed("0001101100011111"),
    signed("0010000101110100"),
    signed("0010001111000101"),
    signed("1101110100010111"),
    signed("0010000101100011"),
    signed("1101011011011110"),
    signed("0010110101010000"),
    signed("1101001010110000"),
    signed("1110011010110011"),
    signed("1110101001001110"),
    signed("0010011110111001"),
    signed("0001111011010101"),
    signed("0001101001000101"),
    signed("1101110111011001"),
    signed("1110010001101000"),
    signed("0010011100110011"),
    signed("1101110011001101"),
    signed("0010010001011111"),
    signed("0001111011000110"),
    signed("0001110010011100"),
    signed("0010001001010000"),
    signed("0010010010111011"),
    signed("1101001010111101"),
    signed("0001111010001011"),
    signed("1110101100101111"),
    signed("0010010000100001"),
    signed("0001110001100010"),
    signed("1101011011101011"),
    signed("1101110010000100"),
    signed("1110001100101101"),
    signed("0001011001000101"),
    signed("0010100001000100"),
    signed("1101101001110010"),
    signed("1110000010001011"),
    signed("0001010101010111"),
    signed("0001110001110111"),
    signed("1101011100111001"));



constant lut_gs2i_data_19 : vector_of_signed16(0 to 63) := 
   (signed("0000000011110001"),
    signed("1111010011001001"),
    signed("1110100011011111"),
    signed("0000111111111101"),
    signed("0001001100111011"),
    signed("0001001001011000"),
    signed("1110000001111110"),
    signed("0001101111011010"),
    signed("0001100110001000"),
    signed("1110111110110011"),
    signed("1110000011010111"),
    signed("1101110001110011"),
    signed("0001111000100101"),
    signed("0011000110001110"),
    signed("0000100101010110"),
    signed("0000110010010011"),
    signed("1110101101100101"),
    signed("0001000011010111"),
    signed("0011000010101011"),
    signed("0000111010011110"),
    signed("1101111111111000"),
    signed("0000111010100001"),
    signed("0001111011000100"),
    signed("0001011001101110"),
    signed("1101001010111100"),
    signed("1101101010111001"),
    signed("0000101010110001"),
    signed("0001111010100000"),
    signed("0010001001111110"),
    signed("0010010110111110"),
    signed("1101110011111001"),
    signed("0001101110111110"),
    signed("1100111001110010"),
    signed("0011001111101100"),
    signed("1100110000010100"),
    signed("1110100101000000"),
    signed("1111010011010110"),
    signed("0010000010000101"),
    signed("0001011000100100"),
    signed("0001010010011011"),
    signed("1110010110011100"),
    signed("1110000000010011"),
    signed("0010010100100010"),
    signed("1110010110011100"),
    signed("0010100000101011"),
    signed("0001110001100000"),
    signed("0001011011110101"),
    signed("0010000010011011"),
    signed("0010101011100111"),
    signed("1100110101110100"),
    signed("0010001101100001"),
    signed("1111001000001101"),
    signed("0010100001111011"),
    signed("0001100010100110"),
    signed("1100111111010010"),
    signed("1101101110011100"),
    signed("1110111100000101"),
    signed("0000100111011101"),
    signed("0010100100101110"),
    signed("1101111111110100"),
    signed("1110101010110010"),
    signed("0000100101010110"),
    signed("0000111100101000"),
    signed("1101000100101110"));



constant lut_gs2i_data_20 : vector_of_signed16(0 to 63) := 
   (signed("0000000100011111"),
    signed("1111110111000111"),
    signed("1111010110100011"),
    signed("0000010100111111"),
    signed("0000110001011100"),
    signed("0000010111010101"),
    signed("1110011000100000"),
    signed("0001101010001100"),
    signed("0000110001110100"),
    signed("1111100000011110"),
    signed("1110110110001010"),
    signed("1101111000011011"),
    signed("0001010100010110"),
    signed("0011011000101110"),
    signed("1111111010101011"),
    signed("0000010111001000"),
    signed("1111001000011111"),
    signed("0000010111000100"),
    signed("0011001000011110"),
    signed("0000001001111111"),
    signed("1110011000110101"),
    signed("0000000110110001"),
    signed("0001111111010100"),
    signed("0000111111000111"),
    signed("1101000010011111"),
    signed("1101011101010110"),
    signed("0000000100010010"),
    signed("0010001101010010"),
    signed("0010001100101010"),
    signed("0010011100000010"),
    signed("1101111000000111"),
    signed("0001001011111110"),
    signed("1100100010010110"),
    signed("0011011100110001"),
    signed("1100100011001111"),
    signed("1110101001001111"),
    signed("1111111101110000"),
    signed("0001010011001001"),
    signed("0000101011011110"),
    signed("0000110111100001"),
    signed("1111000010100101"),
    signed("1101101010110100"),
    signed("0001111010100110"),
    signed("1111000111100000"),
    signed("0010101010000110"),
    signed("0001101001111000"),
    signed("0000111110110010"),
    signed("0001111001110101"),
    signed("0010111110011001"),
    signed("1100101110001111"),
    signed("0010100001110110"),
    signed("1111100010110100"),
    signed("0010110000010101"),
    signed("0001010111100110"),
    signed("1100101101010111"),
    signed("1101101101100101"),
    signed("1111110001111110"),
    signed("1111110101011011"),
    signed("0010011111100111"),
    signed("1110100101111010"),
    signed("1111011110001001"),
    signed("1111110101101111"),
    signed("0000000001100001"),
    signed("1100110110101001"));



constant lut_gs2i_data_21 : vector_of_signed16(0 to 63) := 
   (signed("0000000100011101"),
    signed("0000011000110111"),
    signed("0000001111001001"),
    signed("1111101001100100"),
    signed("0000010010100111"),
    signed("1111100011010100"),
    signed("1110111010111110"),
    signed("0001101000011000"),
    signed("1111110110010010"),
    signed("0000000011001000"),
    signed("1111110011001010"),
    signed("1110000010000000"),
    signed("0000100101100110"),
    signed("0011011111000001"),
    signed("1111010011110101"),
    signed("1111111100111000"),
    signed("1111100111001001"),
    signed("1111101010010001"),
    signed("0011000011001001"),
    signed("1111011001100110"),
    signed("1110111110000110"),
    signed("1111010011110101"),
    signed("0010000011111000"),
    signed("0000011111011101"),
    signed("1101000010101111"),
    signed("1101010011011010"),
    signed("1111100000100011"),
    signed("0010100000100101"),
    signed("0010001101100110"),
    signed("0010011101011101"),
    signed("1101111110111000"),
    signed("0000100000001010"),
    signed("1100010111010001"),
    signed("0011011100101101"),
    signed("1100100011010011"),
    signed("1110100111100110"),
    signed("0000100101100110"),
    signed("0000011000110111"),
    signed("1111111001011010"),
    signed("0000011000110111"),
    signed("1111110110010010"),
    signed("1101010101101110"),
    signed("0001010001111000"),
    signed("0000000000000000"),
    signed("0010101101010011"),
    signed("0001100101010000"),
    signed("0000011100010101"),
    signed("0001110001010001"),
    signed("0011001001010010"),
    signed("1100110011010000"),
    signed("0010110011001100"),
    signed("1111111100111000"),
    signed("0010111001011100"),
    signed("0001010001110101"),
    signed("1100100111001111"),
    signed("1101101111010010"),
    signed("0000101000101110"),
    signed("1111000110111111"),
    signed("0010010100100011"),
    signed("1111010111010010"),
    signed("0000010101101111"),
    signed("1111001010000111"),
    signed("1111000110111111"),
    signed("1100110011010000"));



constant lut_gs2i_data_22 : vector_of_signed16(0 to 63) := 
   (signed("0000000011100111"),
    signed("0000110111100001"),
    signed("0001000101110011"),
    signed("1111000001011000"),
    signed("1111110001000010"),
    signed("1110110010111001"),
    signed("1111100110101100"),
    signed("0001101010001100"),
    signed("1110111011111010"),
    signed("0000100101100111"),
    signed("0000110001100000"),
    signed("1110001011101001"),
    signed("1111110001101001"),
    signed("0011011000101110"),
    signed("1110110011001001"),
    signed("1111100010110100"),
    signed("0000001000111001"),
    signed("1111000000011001"),
    signed("0010110101010001"),
    signed("1110101101111101"),
    signed("1111101100011100"),
    signed("1110100111000011"),
    signed("0010000111101111"),
    signed("1111111011101110"),
    signed("1101001010111001"),
    signed("1101001111100100"),
    signed("1111000000111001"),
    signed("0010101111100100"),
    signed("0010001100101010"),
    signed("0010011010101111"),
    signed("1110000101111000"),
    signed("1111101111111100"),
    signed("1100011001111100"),
    signed("0011010000101011"),
    signed("1100101111010101"),
    signed("1110100000110100"),
    signed("0001001000001111"),
    signed("1111011011011111"),
    signed("1111001000010101"),
    signed("1111110111000111"),
    signed("0000101011001010"),
    signed("1101000110000101"),
    signed("0000011110100100"),
    signed("0000111000100000"),
    signed("0010101010000110"),
    signed("0001100100011100"),
    signed("1111110101111110"),
    signed("0001101010110000"),
    signed("0011001010100000"),
    signed("1101000010110000"),
    signed("0010111101011110"),
    signed("0000010111001000"),
    signed("0010111011001000"),
    signed("0001010010001010"),
    signed("1100101101010111"),
    signed("1101110011000001"),
    signed("0001011010000110"),
    signed("1110100000000011"),
    signed("0010000110111101"),
    signed("0000001110000010"),
    signed("0001001010011010"),
    signed("1110100101110011"),
    signed("1110010011111101"),
    signed("1100111010010101"));



constant lut_gs2i_data_23 : vector_of_signed16(0 to 63) := 
   (signed("0000000010000011"),
    signed("0001010010011011"),
    signed("0001110011001011"),
    signed("1110011111111100"),
    signed("1111001101101001"),
    signed("1110001011100010"),
    signed("0000011000010011"),
    signed("0001101111011010"),
    signed("1110001010111110"),
    signed("0001000110101101"),
    signed("0001101000001111"),
    signed("1110010010100011"),
    signed("1110111110001011"),
    signed("0011000110001110"),
    signed("1110011010011111"),
    signed("1111001000001101"),
    signed("0000101100110111"),
    signed("1110011100100101"),
    signed("0010100001111011"),
    signed("1110001011100010"),
    signed("0000011111111010"),
    signed("1110000101010100"),
    signed("0010001001111110"),
    signed("1111010101001111"),
    signed("1101011001110110"),
    signed("1101010011110101"),
    signed("1110100110010010"),
    signed("0010110101101000"),
    signed("0010001001111110"),
    signed("0010010011101010"),
    signed("1110001010111101"),
    signed("1111000000000011"),
    signed("1100101010111000"),
    signed("0010111010100001"),
    signed("1101000101011111"),
    signed("1110010110000110"),
    signed("0001100011011010"),
    signed("1110100011011111"),
    signed("1110011110000010"),
    signed("1111010011001001"),
    signed("0001011010101010"),
    signed("1101000000101011"),
    signed("1111100101100110"),
    signed("0001101001100100"),
    signed("0010100000101011"),
    signed("0001100111110011"),
    signed("1111001101101001"),
    signed("0001101000000011"),
    signed("0011000000110010"),
    signed("1101011001111001"),
    signed("0010111101001011"),
    signed("0000110010010011"),
    signed("0010110011110001"),
    signed("0001011000111001"),
    signed("1100111111010010"),
    signed("1101111000001001"),
    signed("0010000000001100"),
    signed("1110000011111111"),
    signed("0001111010010001"),
    signed("0001000011111011"),
    signed("0001110101010001"),
    signed("1110001011100101"),
    signed("1101101110110100"),
    signed("1101001010111111"));



constant lut_gs2i_data_24 : vector_of_signed16(0 to 63) := 
   (signed("1111111111111110"),
    signed("0001101001000101"),
    signed("0010010001001001"),
    signed("1110001000001101"),
    signed("1110101001110001"),
    signed("1101110001110110"),
    signed("0001001100000000"),
    signed("0001110111010111"),
    signed("1101101010011110"),
    signed("0001100101001110"),
    signed("0010001111101101"),
    signed("1110010100011111"),
    signed("1110010000011100"),
    signed("0010101000101111"),
    signed("1110001011001011"),
    signed("1110101100101111"),
    signed("0001010001110101"),
    signed("1110000001010000"),
    signed("0010001100010100"),
    signed("1101110110000011"),
    signed("0001010100001000"),
    signed("1101110010011000"),
    signed("0010001010000000"),
    signed("1110101101101101"),
    signed("1101101110010100"),
    signed("1101100001100000"),
    signed("1110010001010011"),
    signed("0010101111001101"),
    signed("0010000101110100"),
    signed("0010001000001101"),
    signed("1110001100010111"),
    signed("1110010100110101"),
    signed("1101001001100001"),
    signed("0010011100011110"),
    signed("1101100011100010"),
    signed("1110001000110110"),
    signed("0001110101010011"),
    signed("1101111000010111"),
    signed("1101111111100010"),
    signed("1110101110001011"),
    signed("0001111111000011"),
    signed("1101001001001000"),
    signed("1110101100000101"),
    signed("0010001100110011"),
    signed("0010010001011111"),
    signed("0001101111001111"),
    signed("1110100101100100"),
    signed("0001101010011000"),
    signed("0010101011101101"),
    signed("1101110101101100"),
    signed("0010101111111110"),
    signed("0001001110110111"),
    signed("0010100010011011"),
    signed("0001100101101011"),
    signed("1101011011101011"),
    signed("1101111101111011"),
    signed("0010010110001110"),
    signed("1101110101010010"),
    signed("0001110001010110"),
    signed("0001110011010011"),
    signed("0010010000101011"),
    signed("1101111101011011"),
    signed("1101011100100000"),
    signed("1101100011101111"));



constant lut_gs2i_data_25 : vector_of_signed16(0 to 63) := 
   (signed("1111111011011101"),
    signed("0001111001000001"),
    signed("0010011001011010"),
    signed("1101111010000111"),
    signed("1110000100111010"),
    signed("1101101011001001"),
    signed("0010000000000001"),
    signed("0001111110111000"),
    signed("1101011100111100"),
    signed("0010000010000110"),
    signed("0010100000011010"),
    signed("1110001110000001"),
    signed("1101101010011001"),
    signed("0010000100010111"),
    signed("1110001000001000"),
    signed("1110010010111011"),
    signed("0001111000011100"),
    signed("1101101101101000"),
    signed("0001110101001110"),
    signed("1101110010001001"),
    signed("0010000010101011"),
    signed("1101101110001100"),
    signed("0010000101100000"),
    signed("1110000100111010"),
    signed("1110001001010000"),
    signed("1101111011000100"),
    signed("1110000100010101"),
    signed("0010011000010001"),
    signed("0001111110011111"),
    signed("0001110110010111"),
    signed("1110001011010111"),
    signed("1101110100000011"),
    signed("1101110001111110"),
    signed("0001111011000110"),
    signed("1110000100111010"),
    signed("1101111000011011"),
    signed("0001111010100011"),
    signed("1101100001110111"),
    signed("1101101110001100"),
    signed("1110000111100100"),
    signed("0010010001110100"),
    signed("1101011111000011"),
    signed("1101110100101000"),
    signed("0010011111110101"),
    signed("0001111111011100"),
    signed("0001110111111000"),
    signed("1101111101111010"),
    signed("0001110100010000"),
    signed("0010001110000010"),
    signed("1110010001001110"),
    signed("0010010010111101"),
    signed("0001101010011011"),
    signed("0010001001010010"),
    signed("0001111001100100"),
    signed("1110000010101001"),
    signed("1110000101110111"),
    signed("0010011011011111"),
    signed("1101110111011101"),
    signed("0001110000010011"),
    signed("0010010101100111"),
    signed("0010011011000110"),
    signed("1101111010000111"),
    signed("1101100001110111"),
    signed("1110000000100100"));



constant lut_gs2i_data_26 : vector_of_signed16(0 to 63) := 
   (signed("1111111001100000"),
    signed("0010001000101011"),
    signed("0010010001001001"),
    signed("1101111101011011"),
    signed("1101100011101111"),
    signed("1101110001110110"),
    signed("0010101101111001"),
    signed("0010001011010111"),
    signed("1101100110101111"),
    signed("0010011001100111"),
    signed("0010011010101100"),
    signed("1110000101110001"),
    signed("1101010001010000"),
    signed("0001011001000101"),
    signed("1110001110111001"),
    signed("1101110101001110"),
    signed("0010011000000100"),
    signed("1101101000100000"),
    signed("0001100101101011"),
    signed("1101111001111111"),
    signed("0010101110010111"),
    signed("1101111111100010"),
    signed("0001111111011011"),
    signed("1101011111110011"),
    signed("1110100010111011"),
    signed("1110011001000010"),
    signed("1101111000100011"),
    signed("0001110111101100"),
    signed("0001110111010011"),
    signed("0001100000111101"),
    signed("1110000101010011"),
    signed("1101011001011000"),
    signed("1110100011111101"),
    signed("0001010110000010"),
    signed("1110101001111110"),
    signed("1101101100111111"),
    signed("0001111001001111"),
    signed("1101100000001111"),
    signed("1101110010011000"),
    signed("1101100111111100"),
    signed("0010010011010000"),
    signed("1110001000100001"),
    signed("1101001001111111"),
    signed("0010011001111100"),
    signed("0001100100110000"),
    signed("0010000111001010"),
    signed("1101011011100111"),
    signed("0001111110010111"),
    signed("0001100110110101"),
    signed("1110110001001001"),
    signed("0001101001111100"),
    signed("0010000110100110"),
    signed("0001100110110001"),
    signed("0010010000000011"),
    signed("1110101110110110"),
    signed("1110001000101101"),
    signed("0010001100110011"),
    signed("1110000111101111"),
    signed("0001110101000100"),
    signed("0010101011000001"),
    signed("0010001100101111"),
    signed("1110001000001101"),
    signed("1101111100000110"),
    signed("1110100110000010"));



constant lut_gs2i_data_27 : vector_of_signed16(0 to 63) := 
   (signed("1111111000011100"),
    signed("0010010001100011"),
    signed("0001110011001011"),
    signed("1110001011100101"),
    signed("1101001010111111"),
    signed("1110001011100010"),
    signed("0011001111101000"),
    signed("0010010100111000"),
    signed("1110001000110111"),
    signed("0010101000010001"),
    signed("0010000010000101"),
    signed("1101110110100110"),
    signed("1101001000010001"),
    signed("0000100111011101"),
    signed("1110011100100110"),
    signed("1101011100000000"),
    signed("0010110101000001"),
    signed("1101101010001100"),
    signed("0001011000111001"),
    signed("1110010011001000"),
    signed("0011001101100010"),
    signed("1110011110000010"),
    signed("0001111011000111"),
    signed("1101000011011001"),
    signed("1111000000111001"),
    signed("1111000000000011"),
    signed("1101110011111001"),
    signed("0001001001011011"),
    signed("0001110011100001"),
    signed("0001001010110100"),
    signed("1101111000101101"),
    signed("1101001100001111"),
    signed("1111011110000000"),
    signed("0000101100110111"),
    signed("1111010011001001"),
    signed("1101100001011011"),
    signed("0001101011000001"),
    signed("1101110000111010"),
    signed("1110000101010100"),
    signed("1101001010111111"),
    signed("0010000101101000"),
    signed("1110111100000101"),
    signed("1100101000110001"),
    signed("0010000010010010"),
    signed("0001001000110100"),
    signed("0010010100111000"),
    signed("1101000011011001"),
    signed("0010001101100001"),
    signed("0000110110010111"),
    signed("1111001101101101"),
    signed("0000111010100001"),
    signed("0010100100000000"),
    signed("0000111010011110"),
    signed("0010100100000001"),
    signed("1111011010101010"),
    signed("1110001100011111"),
    signed("0001101001100100"),
    signed("1110100010000010"),
    signed("0001111100010111"),
    signed("0010110101101000"),
    signed("0001101101101011"),
    signed("1110011111111100"),
    signed("1110100101100101"),
    signed("1111001011100011"));



constant lut_gs2i_data_28 : vector_of_signed16(0 to 63) := 
   (signed("1111111000011110"),
    signed("0010010110000111"),
    signed("0001000101110011"),
    signed("1110100101110011"),
    signed("1100111010010101"),
    signed("1110110010111001"),
    signed("0011100100111011"),
    signed("0010011100010110"),
    signed("1110111100001111"),
    signed("0010101111110111"),
    signed("0001011000000100"),
    signed("1101100101011000"),
    signed("1101001011110101"),
    signed("1111110101011011"),
    signed("1110110010110101"),
    signed("1101000111010111"),
    signed("0011001010100110"),
    signed("1101110010101011"),
    signed("0001010010001010"),
    signed("1110111000101001"),
    signed("0011100000010100"),
    signed("1111001000010101"),
    signed("0001110111001011"),
    signed("1100101111101001"),
    signed("1111100000001010"),
    signed("1111101011000001"),
    signed("1101110011001011"),
    signed("0000010100000111"),
    signed("0001110001011010"),
    signed("0000110001110001"),
    signed("1101101010000000"),
    signed("1101001001110100"),
    signed("0000011000110100"),
    signed("0000000011111110"),
    signed("1111111100000010"),
    signed("1101011001010010"),
    signed("0001010010111011"),
    signed("1110010011101000"),
    signed("1110100111000011"),
    signed("1100110101011010"),
    signed("0001101000010100"),
    signed("1111110110111001"),
    signed("1100010101010101"),
    signed("0001011001110010"),
    signed("0000101010001110"),
    signed("0010100001010010"),
    signed("1100110100100101"),
    signed("0010011100111010"),
    signed("0000000010110001"),
    signed("1111101000111000"),
    signed("0000000110110001"),
    signed("0010111101100101"),
    signed("0000001001111111"),
    signed("0010110100111100"),
    signed("0000000101010101"),
    signed("1110001110100110"),
    signed("0000111000100000"),
    signed("1111000101111111"),
    signed("0010000110101001"),
    signed("0010110100011111"),
    signed("0000111111101110"),
    signed("1111000001011000"),
    signed("1111011011001010"),
    signed("1111110001010110"));



constant lut_gs2i_data_29 : vector_of_signed16(0 to 63) := 
   (signed("1111111001101001"),
    signed("0010010110110111"),
    signed("0000001111001001"),
    signed("1111001010000111"),
    signed("1100110011010000"),
    signed("1111100011010100"),
    signed("0011101100001100"),
    signed("0010100000100101"),
    signed("1111111001011010"),
    signed("0010110000011011"),
    signed("0000100010100101"),
    signed("1101010101101110"),
    signed("1101011000110110"),
    signed("1111000110111111"),
    signed("1111010000101101"),
    signed("1100111001110110"),
    signed("0011010110011101"),
    signed("1101111110111000"),
    signed("0001010001110101"),
    signed("1111100110011100"),
    signed("0011100101100111"),
    signed("1111111001011010"),
    signed("0001110100011001"),
    signed("1100100110011011"),
    signed("0000000000000000"),
    signed("0000010110011100"),
    signed("1101110101001010"),
    signed("1111011101100010"),
    signed("0001110001010001"),
    signed("0000010101101111"),
    signed("1101011100010011"),
    signed("1101010000010010"),
    signed("0001001110110000"),
    signed("1111011101011011"),
    signed("0000100010100101"),
    signed("1101010101101110"),
    signed("0000110010011011"),
    signed("1111000011110111"),
    signed("1111010011110101"),
    signed("1100101001100011"),
    signed("0000111110011101"),
    signed("0000110010011011"),
    signed("1100010000101100"),
    signed("0000100101100110"),
    signed("0000001001101110"),
    signed("0010101010010010"),
    signed("1100110000001000"),
    signed("0010101001011110"),
    signed("1111010000101101"),
    signed("0000000011001000"),
    signed("1111010011110101"),
    signed("0011001111111000"),
    signed("1111011001100110"),
    signed("0011000000000001"),
    signed("0000101100001011"),
    signed("1110001110101111"),
    signed("0000000000000000"),
    signed("1111110000001001"),
    signed("0010010001011011"),
    signed("0010101010010010"),
    signed("0000001000111001"),
    signed("1111101001100100"),
    signed("0000010101101111"),
    signed("0000010101101111"));



constant lut_gs2i_data_30 : vector_of_signed16(0 to 63) := 
   (signed("1111111011110110"),
    signed("0010010100011100"),
    signed("1111010110100011"),
    signed("1111110101101111"),
    signed("1100110110101001"),
    signed("0000010111010101"),
    signed("0011100100111011"),
    signed("0010100000011111"),
    signed("0000110111100100"),
    signed("0010101010011011"),
    signed("1111101000110101"),
    signed("1101001011100001"),
    signed("1101101011001001"),
    signed("1110100000000011"),
    signed("1111110100111010"),
    signed("1100110101110101"),
    signed("0011010110101101"),
    signed("1110001011010100"),
    signed("0001010111100110"),
    signed("0000010111101001"),
    signed("0011011101010101"),
    signed("0000101011011110"),
    signed("0001110011011111"),
    signed("1100101000111111"),
    signed("0000011111110110"),
    signed("0000111110101000"),
    signed("1101111000100010"),
    signed("1110101011111111"),
    signed("0001110011001010"),
    signed("1111110110110010"),
    signed("1101010011000110"),
    signed("1101011101000001"),
    signed("0001111010010010"),
    signed("1110111011001001"),
    signed("0001000100110111"),
    signed("1101010111100111"),
    signed("0000001011011010"),
    signed("1111111011110001"),
    signed("0000000110110001"),
    signed("1100101001010011"),
    signed("0000001100010010"),
    signed("0001100111011100"),
    signed("1100011010110001"),
    signed("1111101100001101"),
    signed("1111101000000100"),
    signed("0010101101110101"),
    signed("1100110110010101"),
    signed("0010110000001000"),
    signed("1110100100111111"),
    signed("0000011101001100"),
    signed("1110100111000011"),
    signed("0011010111100001"),
    signed("1110101101111101"),
    signed("0011000010101110"),
    signed("0001001100110111"),
    signed("1110001100110110"),
    signed("1111000111100000"),
    signed("0000011100100101"),
    signed("0010011001110110"),
    signed("0010011010101000"),
    signed("1111010000011111"),
    signed("0000010100111111"),
    signed("0001001101011000"),
    signed("0000110111001101"));



constant lut_gs2i_data_31 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("0010001111101011"),
    signed("1110100011011111"),
    signed("0000100101010110"),
    signed("1101000100101110"),
    signed("0001001001011000"),
    signed("0011001111101000"),
    signed("0010011011010000"),
    signed("0001101101101111"),
    signed("0010011110100100"),
    signed("1110110010011001"),
    signed("1101001010011000"),
    signed("1101111110001100"),
    signed("1110000011111111"),
    signed("0000011101110000"),
    signed("1100111101001000"),
    signed("0011001010001100"),
    signed("1110010100101001"),
    signed("0001100010100110"),
    signed("0001000111010001"),
    signed("0011001000010101"),
    signed("0001011000100100"),
    signed("0001110100110110"),
    signed("1100110111111011"),
    signed("0000111111000111"),
    signed("0001100000000100"),
    signed("1101111100000011"),
    signed("1110000101010100"),
    signed("0001110110111101"),
    signed("1111010101001111"),
    signed("1101010001101011"),
    signed("1101101100111111"),
    signed("0010010110101001"),
    signed("1110011110101011"),
    signed("0001100001010101"),
    signed("1101011111100011"),
    signed("1111100000001010"),
    signed("0000110101000001"),
    signed("0000111010100001"),
    signed("1100110101110100"),
    signed("1111010110101100"),
    signed("0010001111000110"),
    signed("1100110010011110"),
    signed("1110110100011110"),
    signed("1111000110000110"),
    signed("0010101010001010"),
    signed("1101000110110101"),
    signed("0010101110010001"),
    signed("1110000011111111"),
    signed("0000110111110011"),
    signed("1110000101010100"),
    signed("0011010001110010"),
    signed("1110001011100010"),
    signed("0010111011000101"),
    signed("0001100101100001"),
    signed("1110001001000011"),
    signed("1110010110011100"),
    signed("0001000111010001"),
    signed("0010011101000111"),
    signed("0010001001011010"),
    signed("1110011101111111"),
    signed("0000111111111101"),
    signed("0001111010011111"),
    signed("0001010100100001"));



constant lut_gs2i_data_32 : vector_of_signed16(0 to 63) := 
   (signed("0000000010110111"),
    signed("0010001001011101"),
    signed("1101111100100100"),
    signed("0001010101010111"),
    signed("1101011100111001"),
    signed("0001110100100001"),
    signed("0010101101111001"),
    signed("0010010000010110"),
    signed("0010010100000111"),
    signed("0010001101110000"),
    signed("1110000110000111"),
    signed("1101010100111111"),
    signed("1110001101111010"),
    signed("1101110101010010"),
    signed("0001001001000010"),
    signed("1101010000100101"),
    signed("0010110000110111"),
    signed("1110011000001110"),
    signed("0001110001100010"),
    signed("0001110000110011"),
    signed("0010101000010001"),
    signed("0001111011010101"),
    signed("0001111000100110"),
    signed("1101010010111000"),
    signed("0001011101000101"),
    signed("0001110111110011"),
    signed("1101111110100111"),
    signed("1101101110001100"),
    signed("0001111100010100"),
    signed("1110110001111001"),
    signed("1101011010100111"),
    signed("1101111101001111"),
    signed("0010100000100010"),
    signed("1110001001001011"),
    signed("0001110110110101"),
    signed("1101101101110001"),
    signed("1110110011010000"),
    signed("0001101001101111"),
    signed("0001101001111100"),
    signed("1101001111001001"),
    signed("1110100010100010"),
    signed("0010100011111110"),
    signed("1101010101110110"),
    signed("1110000100100101"),
    signed("1110100100110100"),
    signed("0010011110000110"),
    signed("1101100000101000"),
    signed("0010100010001110"),
    signed("1101110001000110"),
    signed("0001010011010001"),
    signed("1101110010011000"),
    signed("0010111101001011"),
    signed("1101110110000011"),
    signed("0010101000000011"),
    signed("0001110100110101"),
    signed("1110000011101100"),
    signed("1101110011001101"),
    signed("0001101100100110"),
    signed("0010011000111011"),
    signed("0001111010001111"),
    signed("1101111000001010"),
    signed("0001100110111110"),
    signed("0010010110110000"),
    signed("0001101100110100"));



constant lut_gs2i_data_33 : vector_of_signed16(0 to 63) := 
   (signed("0000001001110000"),
    signed("0010000000100101"),
    signed("1101100100100001"),
    signed("0010000000000001"),
    signed("1101111011101001"),
    signed("0010010010111101"),
    signed("0010000000000001"),
    signed("0010000001101101"),
    signed("0010100111011010"),
    signed("0001110110110000"),
    signed("1101100111001011"),
    signed("1101101110101111"),
    signed("1110011001010111"),
    signed("1101110011000111"),
    signed("0001110010000001"),
    signed("1101110001111110"),
    signed("0010001001101011"),
    signed("1110010110101101"),
    signed("0010000000100101"),
    signed("0010001110100111"),
    signed("0001111101010111"),
    signed("0010001101011110"),
    signed("0001111100001110"),
    signed("1101110110010101"),
    signed("0001111011000110"),
    signed("0010000001100011"),
    signed("1101111101010110"),
    signed("1101100111001011"),
    signed("0010000000100101"),
    signed("1110001011111010"),
    signed("1101110001011001"),
    signed("1110001001000110"),
    signed("0010011000110101"),
    signed("1101111000111111"),
    signed("0010000111000001"),
    signed("1110000100010101"),
    signed("1110001001101001"),
    signed("0010010111010011"),
    signed("0010001110100111"),
    signed("1101110001111110"),
    signed("1101110110010101"),
    signed("0010100101001001"),
    signed("1101111111111111"),
    signed("1101100011011001"),
    signed("1110000011001110"),
    signed("0010000111000001"),
    signed("1101111111111111"),
    signed("0010001101101001"),
    signed("1101101100000110"),
    signed("0001101101000101"),
    signed("1101110010100010"),
    signed("0010010111101100"),
    signed("1101101101110011"),
    signed("0010000111100110"),
    signed("0001111100001111"),
    signed("1101111111011011"),
    signed("1101100000001011"),
    signed("0010001011111100"),
    signed("0010001001101011"),
    signed("0001101101101001"),
    signed("1101100001110111"),
    signed("0010000100111100"),
    signed("0010011100000100"),
    signed("0010000001101101"));



constant lut_gs2i_data_34 : vector_of_signed16(0 to 63) := 
   (signed("0000001111001000"),
    signed("0001111000100110"),
    signed("1101100100101000"),
    signed("0010101000101111"),
    signed("1110100101100000"),
    signed("0010100101011001"),
    signed("0001001100000000"),
    signed("0001101000111000"),
    signed("0010100010100111"),
    signed("0001100001000001"),
    signed("1101011111011110"),
    signed("1110010000011100"),
    signed("1110011100011010"),
    signed("1110000100000000"),
    signed("0010011100011010"),
    signed("1110011100111001"),
    signed("0001011001110000"),
    signed("1110001001100000"),
    signed("0010010000100001"),
    signed("0010100101011001"),
    signed("0001001101001110"),
    signed("0010010011010000"),
    signed("0010000101101111"),
    signed("1110100010100010"),
    signed("0010010101011011"),
    signed("0001111110110111"),
    signed("1101111110100111"),
    signed("1101110111011001"),
    signed("0010000101101111"),
    signed("1101100111111100"),
    signed("1110001111001101"),
    signed("1110010001011100"),
    signed("0001111001111001"),
    signed("1101110000101000"),
    signed("0010001111011000"),
    signed("1110011100000101"),
    signed("1101100011100110"),
    signed("0010110011111010"),
    signed("0010101100010000"),
    signed("1110100010100010"),
    signed("1101010010111000"),
    signed("0010001111110001"),
    signed("1110110000010010"),
    signed("1101010000110011"),
    signed("1101101001010111"),
    signed("0001101000001000"),
    signed("1110100101100000"),
    signed("0001101010101101"),
    signed("1101111011111000"),
    signed("0010001010110010"),
    signed("1110000011010000"),
    signed("0001100110000101"),
    signed("1101110110010000"),
    signed("0001100001110100"),
    signed("0001110100110101"),
    signed("1101111010010001"),
    signed("1101100110000100"),
    signed("0010100001000000"),
    signed("0001110001101011"),
    signed("0001100111110010"),
    signed("1101100000011100"),
    signed("0010011110100000"),
    signed("0010001111111010"),
    signed("0010001100011010"));



constant lut_gs2i_data_35 : vector_of_signed16(0 to 63) := 
   (signed("0000010101011001"),
    signed("0001110100110110"),
    signed("1101110110011010"),
    signed("0011000110001110"),
    signed("1111010001010000"),
    signed("0010101110010101"),
    signed("0000011000010011"),
    signed("0001001100111011"),
    signed("0010000100001011"),
    signed("0001000110101101"),
    signed("1101101001010111"),
    signed("1110111110001011"),
    signed("1110010100101001"),
    signed("1110011111111100"),
    signed("0010111110101000"),
    signed("1111001011110000"),
    signed("0000100111001101"),
    signed("1101111000101101"),
    signed("0010100001111011"),
    signed("0010101110010101"),
    signed("0000011101110000"),
    signed("0010000101101000"),
    signed("0010001101100100"),
    signed("1111010110101100"),
    signed("0010101000010001"),
    signed("0001110010010100"),
    signed("1101111100000011"),
    signed("1110010110011100"),
    signed("0010001101100100"),
    signed("1101001010111111"),
    signed("1110111000101111"),
    signed("1110010111111101"),
    signed("0001001101100111"),
    signed("1101110001110011"),
    signed("0010001110001101"),
    signed("1110111010101000"),
    signed("1101000001011000"),
    signed("0011000100110010"),
    signed("0010111011000101"),
    signed("1111010110101100"),
    signed("1100110111111011"),
    signed("0001100100001000"),
    signed("1111100101100110"),
    signed("1101001010011000"),
    signed("1101010010010011"),
    signed("0001000101011000"),
    signed("1111010001010000"),
    signed("0001000010000100"),
    signed("1110011000010101"),
    signed("0010100100000000"),
    signed("1110100000001001"),
    signed("0000101110110100"),
    signed("1110010001000010"),
    signed("0000110010111011"),
    signed("0001100101100001"),
    signed("1101110010011100"),
    signed("1101111101101110"),
    signed("0010101000110101"),
    signed("0001010100010010"),
    signed("0001101011010111"),
    signed("1101110110011010"),
    signed("0010101100001011"),
    signed("0001101101101111"),
    signed("0010010011101010"));



constant lut_gs2i_data_36 : vector_of_signed16(0 to 63) := 
   (signed("0000011101001101"),
    signed("0001110011011111"),
    signed("1110011001101101"),
    signed("0011011000101110"),
    signed("1111111110000100"),
    signed("0010101100111010"),
    signed("1111100110101100"),
    signed("0000101100100001"),
    signed("0001010010110100"),
    signed("0000101010100010"),
    signed("1110000101101110"),
    signed("1111110001101001"),
    signed("1110000110011001"),
    signed("1111000110010011"),
    signed("0011010111111001"),
    signed("1111111100111011"),
    signed("1111110100000010"),
    signed("1101100101000100"),
    signed("0010110000010101"),
    signed("0010101100111010"),
    signed("1111101111111111"),
    signed("0001101000010100"),
    signed("0010010100110001"),
    signed("0000001100010010"),
    signed("0010110100110010"),
    signed("0001011010100001"),
    signed("1101111000100010"),
    signed("1111000010100101"),
    signed("0010010100110001"),
    signed("1100110101011010"),
    signed("1111101000010111"),
    signed("1110011010001100"),
    signed("0000010111001011"),
    signed("1101111000011011"),
    signed("0010000111100101"),
    signed("1111011100011110"),
    signed("1100101000000111"),
    signed("0011001000001010"),
    signed("0010111101110010"),
    signed("0000001100010010"),
    signed("1100101000111111"),
    signed("0000101010010001"),
    signed("0000011001101000"),
    signed("1101010000011100"),
    signed("1101000001111011"),
    signed("0000011110100111"),
    signed("1111111110000100"),
    signed("0000010100101011"),
    signed("1111000000100011"),
    signed("0010111000101001"),
    signed("1111001000000000"),
    signed("1111110100110111"),
    signed("1110111000111101"),
    signed("0000000001000001"),
    signed("0001001100110111"),
    signed("1101101011001111"),
    signed("1110100110001110"),
    signed("0010100110110101"),
    signed("0000110000111000"),
    signed("0001110100101100"),
    signed("1110011110101001"),
    signed("0010110000011100"),
    signed("0000111100100000"),
    signed("0010010101110011"));



constant lut_gs2i_data_37 : vector_of_signed16(0 to 63) := 
   (signed("0000100111010110"),
    signed("0001110100011001"),
    signed("1111001010000111"),
    signed("0011011111000001"),
    signed("0000101000101110"),
    signed("0010100011101101"),
    signed("1110111010111110"),
    signed("0000001000111001"),
    signed("0000010101101111"),
    signed("0000001100110110"),
    signed("1110110001010000"),
    signed("0000100101100110"),
    signed("1101110101001010"),
    signed("1111110011010001"),
    signed("0011100101100111"),
    signed("0000101100001011"),
    signed("1111000100101011"),
    signed("1101010010100110"),
    signed("0010111001011100"),
    signed("0010100011101101"),
    signed("1111000110111111"),
    signed("0000111110011101"),
    signed("0010011001111111"),
    signed("0000111110011101"),
    signed("0010111010001001"),
    signed("0000111001000001"),
    signed("1101110101001010"),
    signed("1111110110010010"),
    signed("0010011001111111"),
    signed("1100101001100011"),
    signed("0000011001100100"),
    signed("1110011000011100"),
    signed("1111011101011011"),
    signed("1110000010000000"),
    signed("0001111110000000"),
    signed("0000000000000000"),
    signed("1100011010011001"),
    signed("0011000000000001"),
    signed("0010110110010100"),
    signed("0000111110011101"),
    signed("1100100110011011"),
    signed("1111101010010001"),
    signed("0001001000001010"),
    signed("1101011111011011"),
    signed("1100111001110110"),
    signed("1111110110010010"),
    signed("0000101000101110"),
    signed("1111100110011100"),
    signed("1111110000001001"),
    signed("0011000110001010"),
    signed("1111110110010010"),
    signed("1110111110000110"),
    signed("1111101001100100"),
    signed("1111010000101101"),
    signed("0000101100001011"),
    signed("1101100110000001"),
    signed("1111011010011010"),
    signed("0010011101011101"),
    signed("0000001001101110"),
    signed("0010000001001000"),
    signed("1111010011110101"),
    signed("0010101100100110"),
    signed("0000000011001000"),
    signed("0010010011101111"));



constant lut_gs2i_data_38 : vector_of_signed16(0 to 63) := 
   (signed("0000110100101001"),
    signed("0001110111001011"),
    signed("0000000001110101"),
    signed("0011011000101110"),
    signed("0001001110000000"),
    signed("0010010110000000"),
    signed("1110011000100000"),
    signed("1111100011101100"),
    signed("1111010101101111"),
    signed("1111101101110100"),
    signed("1111100111001100"),
    signed("0001010100010110"),
    signed("1101100101010101"),
    signed("0000100010010101"),
    signed("0011100101110000"),
    signed("0001010101010001"),
    signed("1110011101011100"),
    signed("1101000101110000"),
    signed("0010111011001000"),
    signed("0010010110000000"),
    signed("1110100101011111"),
    signed("0000001100010010"),
    signed("0010011011111000"),
    signed("0001101000010100"),
    signed("0010110111110001"),
    signed("0000010000000001"),
    signed("1101110011001011"),
    signed("0000101011001010"),
    signed("0010011011111000"),
    signed("1100101001010011"),
    signed("0001000111010111"),
    signed("1110010011100001"),
    signed("1110100111111100"),
    signed("1110001011101001"),
    signed("0001110100010111"),
    signed("0000100011100010"),
    signed("1100011010010000"),
    signed("0010101111100000"),
    signed("0010100111100110"),
    signed("0001101000010100"),
    signed("1100101111101001"),
    signed("1110101101001100"),
    signed("0001101101010000"),
    signed("1101110010101110"),
    signed("1100111011010001"),
    signed("1111001111001000"),
    signed("0001001110000000"),
    signed("1110111011100111"),
    signed("0000100010000001"),
    signed("0011001010001011"),
    signed("0000100101101110"),
    signed("1110010000011010"),
    signed("0000011101011010"),
    signed("1110100110101111"),
    signed("0000000101010101"),
    signed("1101100100001000"),
    signed("0000010011110011"),
    signed("0010001111111100"),
    signed("1111100001011001"),
    signed("0010001101010101"),
    signed("0000001111001011"),
    signed("0010100010101010"),
    signed("1111001001100101"),
    signed("0010001110101100"));



constant lut_gs2i_data_39 : vector_of_signed16(0 to 63) := 
   (signed("0001000101100110"),
    signed("0001111011000111"),
    signed("0000111010100001"),
    signed("0011000110001110"),
    signed("0001101011000001"),
    signed("0010000111010011"),
    signed("1110000001111110"),
    signed("1110111110101111"),
    signed("1110011011111000"),
    signed("1111001101101101"),
    signed("0000100010000000"),
    signed("0001111000100101"),
    signed("1101011011010010"),
    signed("0001001110111000"),
    signed("0011010111001111"),
    signed("0001110100011011"),
    signed("1110000001111110"),
    signed("1101000010110001"),
    signed("0010110011110001"),
    signed("0010000111010011"),
    signed("1110001101101100"),
    signed("1111010110101100"),
    signed("0010011001001010"),
    signed("0010000101101000"),
    signed("0010101101011110"),
    signed("1111100010010000"),
    signed("1101110011111001"),
    signed("0001011010101010"),
    signed("0010011001001010"),
    signed("1100110101110100"),
    signed("0001101100111000"),
    signed("1110001100011111"),
    signed("1101111101111011"),
    signed("1110010010100011"),
    signed("0001101101011101"),
    signed("0001000101011000"),
    signed("1100101000110001"),
    signed("0010011010010100"),
    signed("0010010101000111"),
    signed("0010000101101000"),
    signed("1101000011011001"),
    signed("1101111011110101"),
    signed("0010000101101000"),
    signed("1110000101100000"),
    signed("1101000110110101"),
    signed("1110101011101110"),
    signed("0001101011000001"),
    signed("1110011000010101"),
    signed("0001010000111110"),
    signed("0011000010111000"),
    signed("0001010000111101"),
    signed("1101110000111110"),
    signed("0001001110111000"),
    signed("1110000111011011"),
    signed("1111011010101010"),
    signed("1101100110110110"),
    signed("0001001011100010"),
    signed("0010000001110100"),
    signed("1110111010101000"),
    signed("0010010101110100"),
    signed("0001001001011011"),
    signed("0010010101000111"),
    signed("1110010111110001"),
    signed("0010001000000100"));



constant lut_gs2i_data_40 : vector_of_signed16(0 to 63) := 
   (signed("0001011010010001"),
    signed("0001111111011011"),
    signed("0001101110001001"),
    signed("0010101000101111"),
    signed("0001111101011100"),
    signed("0001111010101101"),
    signed("1101111001000101"),
    signed("1110011100000001"),
    signed("1101110000001111"),
    signed("1110101100111100"),
    signed("0001011100000011"),
    signed("0010001110000101"),
    signed("1101011010110000"),
    signed("0001110100101110"),
    signed("0010111010001101"),
    signed("0010000110110010"),
    signed("1101110100111001"),
    signed("1101001100110111"),
    signed("0010100010011011"),
    signed("0001111010101101"),
    signed("1110000001001001"),
    signed("1110100010100010"),
    signed("0010010000110100"),
    signed("0010010011010000"),
    signed("0010011011100000"),
    signed("1110110010110010"),
    signed("1101111000100011"),
    signed("0001111111000011"),
    signed("0010010000110100"),
    signed("1101001111001001"),
    signed("0010000110000001"),
    signed("1110000100100000"),
    signed("1101100101010100"),
    signed("1110010100011111"),
    signed("0001101011100001"),
    signed("0001100011111011"),
    signed("1101000101110011"),
    signed("0010000100001100"),
    signed("0010000010010011"),
    signed("0010010011010000"),
    signed("1101011111110011"),
    signed("1101011101011001"),
    signed("0010001111000011"),
    signed("1110010011100001"),
    signed("1101011100011011"),
    signed("1110001110010101"),
    signed("0001111101011100"),
    signed("1110000000000100"),
    signed("0001111000011101"),
    signed("0010101111011011"),
    signed("0001110011001100"),
    signed("1101100011011010"),
    signed("0001111000111011"),
    signed("1101110110000111"),
    signed("1110101110110110"),
    signed("1101101111001100"),
    signed("0001111011011011"),
    signed("0001110110010011"),
    signed("1110010111111000"),
    signed("0010010111100000"),
    signed("0001111011111001"),
    signed("0010000110011111"),
    signed("1101110100011111"),
    signed("0010000001010101"));



constant lut_gs2i_data_41 : vector_of_signed16(0 to 63) := 
   (signed("0001110100001011"),
    signed("0010000101100000"),
    signed("0010010101100111"),
    signed("0010000000000001"),
    signed("0010000001100011"),
    signed("0001110100101001"),
    signed("1101111100001100"),
    signed("1101111011010000"),
    signed("1101011010110111"),
    signed("1110001110100100"),
    signed("0010010010011000"),
    signed("0010010000001000"),
    signed("1101100011111110"),
    signed("0010001110100111"),
    signed("0010001110000010"),
    signed("0010001100111001"),
    signed("1101110101001100"),
    signed("1101100011011001"),
    signed("0010000100111100"),
    signed("0001110100101001"),
    signed("1101111110011101"),
    signed("1101110001111110"),
    signed("0010000000000001"),
    signed("0010010001110100"),
    signed("0010000100110000"),
    signed("1110000010101001"),
    signed("1101111111111111"),
    signed("0010010001110100"),
    signed("0010000000000001"),
    signed("1101110110010101"),
    signed("0010001101110111"),
    signed("1101111110110110"),
    signed("1101011111100110"),
    signed("1110010010010111"),
    signed("0001110001111111"),
    signed("0010000000000001"),
    signed("1101101101101000"),
    signed("0001101110001110"),
    signed("0001101111111010"),
    signed("0010010001110100"),
    signed("1110000100111010"),
    signed("1101010100010000"),
    signed("0010001010110100"),
    signed("1110010111101011"),
    signed("1101111000111111"),
    signed("1101110110010101"),
    signed("0010000001100011"),
    signed("1101110011000111"),
    signed("0010010111010011"),
    signed("0010001110000010"),
    signed("0010001010110100"),
    signed("1101100111001011"),
    signed("0010010101100111"),
    signed("1101110110111000"),
    signed("1110000110111111"),
    signed("1101111111111111"),
    signed("0010011100100111"),
    signed("0001101101101001"),
    signed("1101111101010101"),
    signed("0010010010011000"),
    signed("0010011111010001"),
    signed("0001110110111010"),
    signed("1101100110100110"),
    signed("0001111001100100"));



constant lut_gs2i_data_42 : vector_of_signed16(0 to 63) := 
   (signed("0010001101001100"),
    signed("0010001010000000"),
    signed("0010110100011000"),
    signed("0001010101010111"),
    signed("0001111101011100"),
    signed("0001110011101001"),
    signed("1110001101010010"),
    signed("1101100000110001"),
    signed("1101011100000010"),
    signed("1101110001010010"),
    signed("0010111010001101"),
    signed("0010000100111000"),
    signed("1101111110010010"),
    signed("0010100001011110"),
    signed("0001011000010101"),
    signed("0001111111111100"),
    signed("1110000101001001"),
    signed("1110001000100001"),
    signed("0001100011000011"),
    signed("0001110011101001"),
    signed("1110001000001101"),
    signed("1101001111001001"),
    signed("0001101101010010"),
    signed("0001111111000011"),
    signed("0001100111101110"),
    signed("1101010111101111"),
    signed("1110001101100100"),
    signed("0010010011010000"),
    signed("0001101101010010"),
    signed("1110100110010000"),
    signed("0010001001111101"),
    signed("1101110101110011"),
    signed("1101110000010011"),
    signed("1110001001100000"),
    signed("0001111010001111"),
    signed("0010010101111101"),
    signed("1110100011111101"),
    signed("0001100001011111"),
    signed("0001100010101101"),
    signed("0001111111000011"),
    signed("1110101101101101"),
    signed("1101101000001011"),
    signed("0001110110111011"),
    signed("1110010111011101"),
    signed("1110011101010111"),
    signed("1101100111000101"),
    signed("0001111101011100"),
    signed("1101111001001110"),
    signed("0010100101001100"),
    signed("0001100011000111"),
    signed("0010010010110010"),
    signed("1110000010001011"),
    signed("0010101001100110"),
    signed("1110000011010000"),
    signed("1101011111011001"),
    signed("1110010010101110"),
    signed("0010101111001101"),
    signed("0001101011101110"),
    signed("1101100101101001"),
    signed("0001111110110000"),
    signed("0010110111010110"),
    signed("0001101010110110"),
    signed("1101101101011100"),
    signed("0001110100011001"));



constant lut_gs2i_data_43 : vector_of_signed16(0 to 63) := 
   (signed("0010100101000100"),
    signed("0010001001111110"),
    signed("0011000010101011"),
    signed("0000100101010110"),
    signed("0001101011000001"),
    signed("0001110101000011"),
    signed("1110101100111100"),
    signed("1101010000011011"),
    signed("1101110000111010"),
    signed("1101010100011001"),
    signed("0011010111001111"),
    signed("0001100111011110"),
    signed("1110100010000001"),
    signed("0010100110101110"),
    signed("0000011111111010"),
    signed("0001100111101011"),
    signed("1110100101010110"),
    signed("1110111100000101"),
    signed("0000111000010111"),
    signed("0001110101000011"),
    signed("1110011111111100"),
    signed("1100110101110100"),
    signed("0001010010011011"),
    signed("0001011010101010"),
    signed("0001000011010111"),
    signed("1100110111101011"),
    signed("1110100100001011"),
    signed("0010000101101000"),
    signed("0001010010011011"),
    signed("1111011000110011"),
    signed("0001110100011110"),
    signed("1101110000100010"),
    signed("1110010111110001"),
    signed("1101111000101101"),
    signed("0010001001011010"),
    signed("0010100010100100"),
    signed("1111011110000000"),
    signed("0001011000111001"),
    signed("0001011110010110"),
    signed("0001011010101010"),
    signed("1111010101001111"),
    signed("1110010000001011"),
    signed("0001010011000100"),
    signed("1110001101000110"),
    signed("1111001001101001"),
    signed("1101100010111001"),
    signed("0001101011000001"),
    signed("1110001011100101"),
    signed("0010101000110101"),
    signed("0000110100010000"),
    signed("0010000111101111"),
    signed("1110101010110010"),
    signed("0010101110010101"),
    signed("1110100000001001"),
    signed("1101000001011000"),
    signed("1110101101100101"),
    signed("0010110101101000"),
    signed("0001110010111101"),
    signed("1101010111111100"),
    signed("0001100011011011"),
    signed("0010111101001111"),
    signed("0001100101111100"),
    signed("1110000101100001"),
    signed("0001110100110110"));



constant lut_gs2i_data_44 : vector_of_signed16(0 to 63) := 
   (signed("0010111001000110"),
    signed("0010000111101111"),
    signed("0011000011100010"),
    signed("1111110101101111"),
    signed("0001001110000000"),
    signed("0001111010001000"),
    signed("1111010101101011"),
    signed("1101001000100100"),
    signed("1110011000100100"),
    signed("1100111100101011"),
    signed("0011100101110000"),
    signed("0000111101110000"),
    signed("1111001110100111"),
    signed("0010100010001110"),
    signed("1111100111100001"),
    signed("0001000100011001"),
    signed("1111001111111011"),
    signed("1111110110111001"),
    signed("0000001010010011"),
    signed("0001111010001000"),
    signed("1111000001011000"),
    signed("1100101001010011"),
    signed("0000110010100101"),
    signed("0000101011001010"),
    signed("0000011100000000"),
    signed("1100100010101011"),
    signed("1111000001001110"),
    signed("0001101000010100"),
    signed("0000110010100101"),
    signed("0000001011111110"),
    signed("0001010010000011"),
    signed("1101101101010001"),
    signed("1111001110100000"),
    signed("1101100101000100"),
    signed("0010011010101000"),
    signed("0010101000000101"),
    signed("0000011000110100"),
    signed("0001010111000110"),
    signed("0001100000011000"),
    signed("0000101011001010"),
    signed("1111111011101110"),
    signed("1111001000110000"),
    signed("0000100101011001"),
    signed("1101111101011010"),
    signed("1111111000010100"),
    signed("1101100110001010"),
    signed("0001001110000000"),
    signed("1110101010101111"),
    signed("0010100001111001"),
    signed("0000000011000101"),
    signed("0001101100111100"),
    signed("1111011110001001"),
    signed("0010100111111110"),
    signed("1111001000000000"),
    signed("1100101101000010"),
    signed("1111001101011011"),
    signed("0010101111100100"),
    signed("0001111111011000"),
    signed("1101010001110111"),
    signed("0000111111100111"),
    signed("0010110101010100"),
    signed("0001100110001001"),
    signed("1110101101101100"),
    signed("0001111000011010"));



constant lut_gs2i_data_45 : vector_of_signed16(0 to 63) := 
   (signed("0011000110011001"),
    signed("0010000011111000"),
    signed("0010111001011100"),
    signed("1111001010000111"),
    signed("0000101000101110"),
    signed("0010000001001000"),
    signed("0000000011001000"),
    signed("1101001000111111"),
    signed("1111001101100101"),
    signed("1100101101000000"),
    signed("0011100101100111"),
    signed("0000001100110110"),
    signed("0000000000000000"),
    signed("0010010110110111"),
    signed("1110110100011000"),
    signed("0000011001100100"),
    signed("0000000000000000"),
    signed("0000110010011011"),
    signed("1111011100101110"),
    signed("0010000001001000"),
    signed("1111101001100100"),
    signed("1100101001100011"),
    signed("0000001111001001"),
    signed("1111110110010010"),
    signed("1111110011111111"),
    signed("1100011010011001"),
    signed("1111100011101011"),
    signed("0000111110011101"),
    signed("0000001111001001"),
    signed("0000111011010101"),
    signed("0000100110011010"),
    signed("1101101100001010"),
    signed("0000001100110110"),
    signed("1101010010100110"),
    signed("0010101010010010"),
    signed("0010100111001010"),
    signed("0001001110110000"),
    signed("0001011011100010"),
    signed("0001100111100100"),
    signed("1111110110010010"),
    signed("0000011111011101"),
    signed("0000001001101110"),
    signed("1111110011001010"),
    signed("1101101100010001"),
    signed("0000100101100110"),
    signed("1101101110100101"),
    signed("0000101000101110"),
    signed("1111010011110101"),
    signed("0010010011101111"),
    signed("1111010011110101"),
    signed("0001000101000010"),
    signed("0000010101101111"),
    signed("0010011001111111"),
    signed("1111110110010010"),
    signed("1100100100000111"),
    signed("1111110000110111"),
    signed("0010100000100101"),
    signed("0010001101111110"),
    signed("1101010010100110"),
    signed("0000010101101111"),
    signed("0010100011101101"),
    signed("0001101010101100"),
    signed("1111100000100011"),
    signed("0001111110000111"));



constant lut_gs2i_data_46 : vector_of_signed16(0 to 63) := 
   (signed("0011001010001111"),
    signed("0001111111010100"),
    signed("0010100111111011"),
    signed("1110100101110011"),
    signed("1111111110000100"),
    signed("0010000111111001"),
    signed("0000110000011010"),
    signed("1101010000111110"),
    signed("0000001001000111"),
    signed("1100101000001010"),
    signed("0011010111111001"),
    signed("1111011010100111"),
    signed("0000110001011001"),
    signed("0010001000010110"),
    signed("1110001011011111"),
    signed("1111101011010101"),
    signed("0000110000000101"),
    signed("0001100111011100"),
    signed("1110110011101101"),
    signed("0010000111111001"),
    signed("0000010100111111"),
    signed("1100110101011010"),
    signed("1111101001110001"),
    signed("1111000010100101"),
    signed("1111001101101111"),
    signed("1100011111101100"),
    signed("0000001010000010"),
    signed("0000001100010010"),
    signed("1111101001110001"),
    signed("0001100010100100"),
    signed("1111110110000001"),
    signed("1101101101010001"),
    signed("0001001001110110"),
    signed("1101000101110000"),
    signed("0010110100011111"),
    signed("0010100000111110"),
    signed("0001111010010010"),
    signed("0001100100111100"),
    signed("0001110001111010"),
    signed("1111000010100101"),
    signed("0000111111000111"),
    signed("0001001001100010"),
    signed("1111000010010000"),
    signed("1101011110000111"),
    signed("0001001101101011"),
    signed("1101111001010111"),
    signed("1111111110000100"),
    signed("0000000011000101"),
    signed("0010000010100110"),
    signed("1110101010101111"),
    signed("0000010011111000"),
    signed("0001001010011010"),
    signed("0010001000101010"),
    signed("0000100101101110"),
    signed("1100100111100111"),
    signed("0000010110001111"),
    signed("0010001101010010"),
    signed("0010011010111111"),
    signed("1101011000111110"),
    signed("1111101000111100"),
    signed("0010001101100110"),
    signed("0001110010001111"),
    signed("0000010111100000"),
    signed("0010000100100001"));



constant lut_gs2i_data_47 : vector_of_signed16(0 to 63) := 
   (signed("0011000010101000"),
    signed("0001111011000100"),
    signed("0010010011000001"),
    signed("1110001011100101"),
    signed("1111010001010000"),
    signed("0010001100000111"),
    signed("0001011000100100"),
    signed("1101011111010101"),
    signed("0001000011111011"),
    signed("1100110000010100"),
    signed("0010111110101000"),
    signed("1110101100111100"),
    signed("0001011101111111"),
    signed("0001111010100000"),
    signed("1101110000111110"),
    signed("1110111101111100"),
    signed("0001011010101010"),
    signed("0010001111000110"),
    signed("1110010011001000"),
    signed("0010001100000111"),
    signed("0000111111111101"),
    signed("1101001010111111"),
    signed("1111000100001111"),
    signed("1110010110011100"),
    signed("1110101011011111"),
    signed("1100110010011110"),
    signed("0000110010010111"),
    signed("1111010110101100"),
    signed("1111000100001111"),
    signed("0001111110000010"),
    signed("1111000101100010"),
    signed("1101110000100010"),
    signed("0001111100101001"),
    signed("1101000010110001"),
    signed("0010110101101000"),
    signed("0010010110111110"),
    signed("0010010110101001"),
    signed("0001110001100000"),
    signed("0001111101001110"),
    signed("1110010110011100"),
    signed("0001011001101110"),
    signed("0001111110101111"),
    signed("1110011000100010"),
    signed("1101010111001011"),
    signed("0001101101000111"),
    signed("1110000011101001"),
    signed("1111010001010000"),
    signed("0000110100010000"),
    signed("0001110010111010"),
    signed("1110001011100101"),
    signed("1111011110000000"),
    signed("0001110101010001"),
    signed("0001111000011001"),
    signed("0001010000111101"),
    signed("1100110111101011"),
    signed("0000111011110001"),
    signed("0001111010100000"),
    signed("0010100010100111"),
    signed("1101100011100010"),
    signed("1110111100101001"),
    signed("0001111000011001"),
    signed("0001111011000111"),
    signed("0001001011100001"),
    signed("0010001010000001"));



constant lut_gs2i_data_48 : vector_of_signed16(0 to 63) := 
   (signed("0010101110100011"),
    signed("0001111000000100"),
    signed("0001111110100100"),
    signed("1101111101011011"),
    signed("1110100101100000"),
    signed("0010001011101001"),
    signed("0001110111001000"),
    signed("1101110010101110"),
    signed("0001110111011111"),
    signed("1101000110100011"),
    signed("0010011100011010"),
    signed("1110001001000101"),
    signed("0010000001101110"),
    signed("0001110000101011"),
    signed("1101100111100110"),
    signed("1110010101010011"),
    signed("0001111010110111"),
    signed("0010100011111110"),
    signed("1101111110001011"),
    signed("0010001011101001"),
    signed("0001100110111110"),
    signed("1101100111111100"),
    signed("1110100000011011"),
    signed("1101110111011001"),
    signed("1110001111000000"),
    signed("1101010001101001"),
    signed("0001011010011100"),
    signed("1110100010100010"),
    signed("1110100000011011"),
    signed("0010001011000111"),
    signed("1110011001001111"),
    signed("1101110101110011"),
    signed("0010011101101010"),
    signed("1101001100110111"),
    signed("0010101011000001"),
    signed("0010001010111001"),
    signed("0010100000100010"),
    signed("0001111111010010"),
    signed("0010000111010110"),
    signed("1101110111011001"),
    signed("0001101110101101"),
    signed("0010100001011001"),
    signed("1101111011001000"),
    signed("1101011010110100"),
    signed("0010000001001010"),
    signed("1110001010111100"),
    signed("1110100101100000"),
    signed("0001100011000111"),
    signed("0001101000100011"),
    signed("1101111001001110"),
    signed("1110101000001001"),
    signed("0010010000101011"),
    signed("0001101100111101"),
    signed("0001110011001100"),
    signed("1101010011100011"),
    signed("0001011111100101"),
    signed("0001101100011111"),
    signed("0010100001100010"),
    signed("1101110000101110"),
    signed("1110010100000110"),
    signed("0001101000110000"),
    signed("0010000011101000"),
    signed("0001110110001010"),
    signed("0010001101001011"));



constant lut_gs2i_data_49 : vector_of_signed16(0 to 63) := 
   (signed("0010001100001001"),
    signed("0001110100110101"),
    signed("0001101111111010"),
    signed("1101111110011101"),
    signed("1101111111111111"),
    signed("0010000010101011"),
    signed("0010000110011110"),
    signed("1110001011111010"),
    signed("0010011100100111"),
    signed("1101101000010100"),
    signed("0001110110010111"),
    signed("1101110101001100"),
    signed("0010010111101100"),
    signed("0001101111010101"),
    signed("1101110010100010"),
    signed("1101110010010111"),
    signed("0010001111001010"),
    signed("0010100000110011"),
    signed("1101111001001001"),
    signed("0010000010101011"),
    signed("0010001001010010"),
    signed("1110000111100100"),
    signed("1110000010010000"),
    signed("1101101011100010"),
    signed("1101111011101001"),
    signed("1101111101010101"),
    signed("0001111101110000"),
    signed("1101110001111110"),
    signed("1101111101111010"),
    signed("0010001010110100"),
    signed("1101110110101110"),
    signed("1101111110110110"),
    signed("0010100101101110"),
    signed("1101100111101111"),
    signed("0010010101100111"),
    signed("0001111100001110"),
    signed("0010011000110101"),
    signed("0010001110100101"),
    signed("0010010000110110"),
    signed("1101100111001011"),
    signed("0010000000000001"),
    signed("0010101110011010"),
    signed("1101101011100010"),
    signed("1101101000101101"),
    signed("0010000101111001"),
    signed("1110001111101101"),
    signed("1101111011101001"),
    signed("0010001001101011"),
    signed("0001101000010101"),
    signed("1101110011000111"),
    signed("1101110100101000"),
    signed("0010010110110000"),
    signed("0001100110101001"),
    signed("0010001010110100"),
    signed("1101111011101001"),
    signed("0001111101110000"),
    signed("0001101000010101"),
    signed("0010010011010110"),
    signed("1101111100110001"),
    signed("1101101111111001"),
    signed("0001100011111111"),
    signed("0010001100100000"),
    signed("0010010100011110"),
    signed("0010001111001010"));



constant lut_gs2i_data_50 : vector_of_signed16(0 to 63) := 
   (signed("0001100001110110"),
    signed("0001110100010101"),
    signed("0001100110011100"),
    signed("1110001011111011"),
    signed("1101100000101000"),
    signed("0001110110110101"),
    signed("0010001011000111"),
    signed("1110100111000111"),
    signed("0010110011001001"),
    signed("1110010110001101"),
    signed("0001001100110000"),
    signed("1101110000111101"),
    signed("0010100001100010"),
    signed("0001110000101011"),
    signed("1110001110000010"),
    signed("1101011101110010"),
    signed("0010001110110110"),
    signed("0010001100000011"),
    signed("1101111110001011"),
    signed("0001110110110101"),
    signed("0010100010001110"),
    signed("1110101110001011"),
    signed("1101101000101100"),
    signed("1101110001111011"),
    signed("1101101111001100"),
    signed("1110101011111000"),
    signed("0010100000101011"),
    signed("1101001111001001"),
    signed("1101100100111110"),
    signed("0001111010110111"),
    signed("1101011101100101"),
    signed("1110000100100000"),
    signed("0010011001101110"),
    signed("1110001100001111"),
    signed("0001110011010011"),
    signed("0001101111001111"),
    signed("0001111001111001"),
    signed("0010010111001101"),
    signed("0010010010001000"),
    signed("1101101110001100"),
    signed("0010001011001011"),
    signed("0010011101011101"),
    signed("1101101110001100"),
    signed("1110000111100011"),
    signed("0001111101011100"),
    signed("1110001110101010"),
    signed("1101011100111001"),
    signed("0010101011101101"),
    signed("0001101100011111"),
    signed("1110000000000100"),
    signed("1101001101111011"),
    signed("0010001001000000"),
    signed("0001101100111101"),
    signed("0010010010110010"),
    signed("1110101010101001"),
    signed("0010010111010100"),
    signed("0001101000100011"),
    signed("0001111110000000"),
    signed("1110001000110110"),
    signed("1101011000101001"),
    signed("0001101000100011"),
    signed("0010010010001000"),
    signed("0010100000100010"),
    signed("0010001100111110"));



constant lut_gs2i_data_51 : vector_of_signed16(0 to 63) := 
   (signed("0000110000110111"),
    signed("0001111000111101"),
    signed("0001100000011100"),
    signed("1110100010000010"),
    signed("1101000110110101"),
    signed("0001100001010101"),
    signed("0001111110000010"),
    signed("1111000000111001"),
    signed("0010111101001111"),
    signed("1111001111000110"),
    signed("0000011111110110"),
    signed("1101111010011000"),
    signed("0010100010100111"),
    signed("0001111010100000"),
    signed("1110110100011111"),
    signed("1101010001101111"),
    signed("0010000000001000"),
    signed("0001100010000001"),
    signed("1110010011001000"),
    signed("0001100001010101"),
    signed("0010101110010001"),
    signed("1111010011001001"),
    signed("1101010010100010"),
    signed("1110000111011011"),
    signed("1101100110110110"),
    signed("1111100000000110"),
    signed("0010111010100001"),
    signed("1100110101110100"),
    signed("1101010000011011"),
    signed("0001011010101010"),
    signed("1101001100001111"),
    signed("1110001100011111"),
    signed("0001110101000010"),
    signed("1110111110001011"),
    signed("0001000011111011"),
    signed("0001100111110011"),
    signed("0001001101100111"),
    signed("0010011110100101"),
    signed("0010010001100100"),
    signed("1110000101010100"),
    signed("0010001110001101"),
    signed("0001110111001001"),
    signed("1110000101010100"),
    signed("1110101111000010"),
    signed("0001101011000001"),
    signed("1110000101101111"),
    signed("1101000100101110"),
    signed("0011000000110010"),
    signed("0001111010100000"),
    signed("1110011000010101"),
    signed("1100110000011000"),
    signed("0001101011100101"),
    signed("0001111000011001"),
    signed("0010000111101111"),
    signed("1111011010101010"),
    signed("0010101101011110"),
    signed("0001110010111010"),
    signed("0001011011111000"),
    signed("1110010110000110"),
    signed("1101001000110101"),
    signed("0001110010111010"),
    signed("0010010001100100"),
    signed("0010010110101001"),
    signed("0010000100100001"));



constant lut_gs2i_data_52 : vector_of_signed16(0 to 63) := 
   (signed("1111111101011010"),
    signed("0001111111101001"),
    signed("0001100000000100"),
    signed("1111000001000011"),
    signed("1100110110010101"),
    signed("0001000100110111"),
    signed("0001100010100100"),
    signed("1111011011001110"),
    signed("0010111010010000"),
    signed("0000001011011110"),
    signed("1111110100100110"),
    signed("1110010010110000"),
    signed("0010011010111111"),
    signed("0010001000010110"),
    signed("1111100011100101"),
    signed("1101001111111000"),
    signed("0001100010010000"),
    signed("0000101010100110"),
    signed("1110110011101101"),
    signed("0001000100110111"),
    signed("0010110000001000"),
    signed("1111110111000111"),
    signed("1101000011010100"),
    signed("1110101011101010"),
    signed("1101100100001000"),
    signed("0000010011100100"),
    signed("0011001011101111"),
    signed("1100101001010011"),
    signed("1101000011101000"),
    signed("0000110000000101"),
    signed("1101000100111000"),
    signed("1110010011100001"),
    signed("0000111111001010"),
    signed("1111110110100101"),
    signed("0000001110000010"),
    signed("0001100100011100"),
    signed("0000010111001011"),
    signed("0010100001110010"),
    signed("0010001101011111"),
    signed("1110101011111111"),
    signed("0010001100100000"),
    signed("0000111110110110"),
    signed("1110101011111111"),
    signed("1111011101111111"),
    signed("0001001110000000"),
    signed("1101111001000011"),
    signed("1100110110101001"),
    signed("0011001010100000"),
    signed("0010001101010010"),
    signed("1110111011100111"),
    signed("1100100000000001"),
    signed("0001000000000010"),
    signed("0010001000101010"),
    signed("0001101100111100"),
    signed("0000001010010001"),
    signed("0010111100101100"),
    signed("0010000010100110"),
    signed("0000110001101101"),
    signed("1110100000110100"),
    signed("1101000010110011"),
    signed("0010000010100110"),
    signed("0010001101011111"),
    signed("0001111010010010"),
    signed("0001111001100000"));



constant lut_gs2i_data_53 : vector_of_signed16(0 to 63) := 
   (signed("1111001100010000"),
    signed("0010000111000000"),
    signed("0001100100011100"),
    signed("1111100110011100"),
    signed("1100110000001000"),
    signed("0000100010100101"),
    signed("0000111011010101"),
    signed("1111110110010010"),
    signed("0010101101011010"),
    signed("0001000101000010"),
    signed("1111001101100101"),
    signed("1110110111110110"),
    signed("0010001101111110"),
    signed("0010010110110111"),
    signed("0000010101101111"),
    signed("1101010110100010"),
    signed("0000111000001101"),
    signed("1111101101011001"),
    signed("1111011100101110"),
    signed("0000100010100101"),
    signed("0010101001011110"),
    signed("0000011000110111"),
    signed("1100111100001010"),
    signed("1111011010011010"),
    signed("1101100110000001"),
    signed("0001000001111010"),
    signed("0011010011000000"),
    signed("1100101001100011"),
    signed("1100111111010010"),
    signed("0000000000000000"),
    signed("1101000110100100"),
    signed("1110011000011100"),
    signed("0000000000000000"),
    signed("0000101111010011"),
    signed("1111010111010010"),
    signed("0001100101010000"),
    signed("1111011101011011"),
    signed("0010100000100101"),
    signed("0010000111000000"),
    signed("1111011101100010"),
    signed("0010000111101110"),
    signed("1111111100111000"),
    signed("1111011101100010"),
    signed("0000001111110111"),
    signed("0000101000101110"),
    signed("1101101011011101"),
    signed("1100110011010000"),
    signed("0011001001010010"),
    signed("0010100000100101"),
    signed("1111100110011100"),
    signed("1100011101100001"),
    signed("0000001100000001"),
    signed("0010011001111111"),
    signed("0001000101000010"),
    signed("0000110101111001"),
    signed("0011000011110110"),
    signed("0010010011101111"),
    signed("0000000011001000"),
    signed("1110100111100110"),
    signed("1101000101110111"),
    signed("0010010011101111"),
    signed("0010000111000000"),
    signed("0001001110110000"),
    signed("0001101110001001"));



constant lut_gs2i_data_54 : vector_of_signed16(0 to 63) := 
   (signed("1110100010001111"),
    signed("0010001101011111"),
    signed("0001101100001010"),
    signed("0000001111001111"),
    signed("1100110100100101"),
    signed("1111111100000010"),
    signed("0000001011111110"),
    signed("0000010010100000"),
    signed("0010011010111100"),
    signed("0001110101010110"),
    signed("1110101101000101"),
    signed("1111100110011000"),
    signed("0001111111011000"),
    signed("0010100010001110"),
    signed("0001000100111110"),
    signed("1101100011000110"),
    signed("0000000110001110"),
    signed("1110110010111100"),
    signed("0000001010010011"),
    signed("1111111100000010"),
    signed("0010011100111010"),
    signed("0000110111100001"),
    signed("1100111101111000"),
    signed("0000001110010111"),
    signed("1101101011001111"),
    signed("0001100111001011"),
    signed("0011001111011011"),
    signed("1100110101011010"),
    signed("1101000011101000"),
    signed("1111001111111011"),
    signed("1101001111101011"),
    signed("1110011010001100"),
    signed("1111000000110110"),
    signed("0001100001101100"),
    signed("1110100101111010"),
    signed("0001101001111000"),
    signed("1110100111111100"),
    signed("0010011011000011"),
    signed("0001111111101001"),
    signed("0000010100000111"),
    signed("0010000001101101"),
    signed("1110111011000110"),
    signed("0000010100000111"),
    signed("0000111111011101"),
    signed("1111111110000100"),
    signed("1101100000011001"),
    signed("1100111010010101"),
    signed("0010111110011001"),
    signed("0010101111100100"),
    signed("0000010100101011"),
    signed("1100101000011011"),
    signed("1111010110001111"),
    signed("0010100111111110"),
    signed("0000010011111000"),
    signed("0001011010001101"),
    signed("0011000010001000"),
    signed("0010100001111001"),
    signed("1111010100011000"),
    signed("1110101001001111"),
    signed("1101010000101010"),
    signed("0010100001111001"),
    signed("0001111111101001"),
    signed("0000011000110100"),
    signed("0001100101000000"));



constant lut_gs2i_data_55 : vector_of_signed16(0 to 63) := 
   (signed("1110000011101001"),
    signed("0010010001100100"),
    signed("0001110101100111"),
    signed("0000111000010111"),
    signed("1101000011011001"),
    signed("1111010011001001"),
    signed("1111011000110011"),
    signed("0000110000001101"),
    signed("0010000111010011"),
    signed("0010010110101001"),
    signed("1110010100111111"),
    signed("0000011010011010"),
    signed("0001110010111101"),
    signed("0010100110101110"),
    signed("0001101011100101"),
    signed("1101110010011111"),
    signed("1111010001001100"),
    signed("1110000011011011"),
    signed("0000111000010111"),
    signed("1111010011001001"),
    signed("0010001101100001"),
    signed("0001010010011011"),
    signed("1101001000110101"),
    signed("0001000001110101"),
    signed("1101110010011100"),
    signed("0010000000001000"),
    signed("0011000000110010"),
    signed("1101001010111111"),
    signed("1101010000011011"),
    signed("1110100101010110"),
    signed("1101011110000101"),
    signed("1110010111111101"),
    signed("1110001010111110"),
    signed("0010000111011111"),
    signed("1101111111110100"),
    signed("0001110001100000"),
    signed("1101111101111011"),
    signed("0010010001100011"),
    signed("0001111000111101"),
    signed("0001001001011011"),
    signed("0001111100010111"),
    signed("1110000011010111"),
    signed("0001001001011011"),
    signed("0001100111101011"),
    signed("1111010001010000"),
    signed("1101011011010010"),
    signed("1101001010111111"),
    signed("0010101011100111"),
    signed("0010110101101000"),
    signed("0001000010000100"),
    signed("1100111111010010"),
    signed("1110100101100101"),
    signed("0010101110010101"),
    signed("1111011110000000"),
    signed("0001110100011011"),
    signed("0010110111001011"),
    signed("0010101000110101"),
    signed("1110101001101000"),
    signed("1110100101000000"),
    signed("1101100001011100"),
    signed("0010101000110101"),
    signed("0001111000111101"),
    signed("1111011110000000"),
    signed("0001100000011100"));



constant lut_gs2i_data_56 : vector_of_signed16(0 to 63) := 
   (signed("1101110011101000"),
    signed("0010010010001000"),
    signed("0001111111001110"),
    signed("0001011110110110"),
    signed("1101011011100111"),
    signed("1110101001111110"),
    signed("1110100110010000"),
    signed("0001001111010101"),
    signed("0001110110100000"),
    signed("0010100100101110"),
    signed("1110000110110001"),
    signed("0001001111101110"),
    signed("0001101011101110"),
    signed("0010100001011110"),
    signed("0010000100110100"),
    signed("1110000001101001"),
    signed("1110011110001000"),
    signed("1101100101100001"),
    signed("0001100011000011"),
    signed("1110101001111110"),
    signed("0001111110010111"),
    signed("0001101001000101"),
    signed("1101011100110101"),
    signed("0001101111100100"),
    signed("1101111010010001"),
    signed("0010001010101010"),
    signed("0010100111100000"),
    signed("1101100111111100"),
    signed("1101100100111110"),
    signed("1110000101001001"),
    signed("1101101111011111"),
    signed("1110010001011100"),
    signed("1101100110010010"),
    signed("0010011011110101"),
    signed("1101101001110010"),
    signed("0001111011000110"),
    signed("1101100101010100"),
    signed("0010000100011111"),
    signed("0001110100010101"),
    signed("0001110111101100"),
    signed("0001111001010001"),
    signed("1101011110001001"),
    signed("0001110111101100"),
    signed("0010000100001000"),
    signed("1110100101100000"),
    signed("1101011110111100"),
    signed("1101100011101111"),
    signed("0010010010111011"),
    signed("0010101111001101"),
    signed("0001101010101101"),
    signed("1101011111110111"),
    signed("1110000000010010"),
    signed("0010101001100110"),
    signed("1110101000001001"),
    signed("0010000010100101"),
    signed("0010100011001011"),
    signed("0010100101001100"),
    signed("1110000110011010"),
    signed("1110011010110011"),
    signed("1101110110011100"),
    signed("0010100101001100"),
    signed("0001110100010101"),
    signed("1110100011111101"),
    signed("0001100010001111"));



constant lut_gs2i_data_57 : vector_of_signed16(0 to 63) := 
   (signed("1101110001101100"),
    signed("0010010000110110"),
    signed("0010000101100000"),
    signed("0010000010010010"),
    signed("1101111001100100"),
    signed("1110000000100100"),
    signed("1101110110010101"),
    signed("0001101101000101"),
    signed("0001101001010011"),
    signed("0010011111110101"),
    signed("1110000101011101"),
    signed("0010000100010111"),
    signed("0001101101101001"),
    signed("0010001110100111"),
    signed("0010001111101111"),
    signed("1110001011110000"),
    signed("1101110011101011"),
    signed("1101011011010000"),
    signed("0010000100111100"),
    signed("1110000000100100"),
    signed("0001101111111010"),
    signed("0001111001000001"),
    signed("1101111011010000"),
    signed("0010010001010001"),
    signed("1101111111011011"),
    signed("0010001000001010"),
    signed("0010000111000001"),
    signed("1110000111100100"),
    signed("1110000010010000"),
    signed("1101110101001100"),
    signed("1110000011110010"),
    signed("1110000100110000"),
    signed("1101011010010010"),
    signed("0010011001110011"),
    signed("1101101000110111"),
    signed("0010000111100101"),
    signed("1101011111100110"),
    signed("0001110010000001"),
    signed("0001110100110101"),
    signed("0010011100100111"),
    signed("0001110111010011"),
    signed("1101010011010010"),
    signed("0010011100100111"),
    signed("0010010011111010"),
    signed("1101111011101001"),
    signed("1101101111010100"),
    signed("1110000000100100"),
    signed("0001111000011100"),
    signed("0010011000010001"),
    signed("0010001101101001"),
    signed("1110000101010011"),
    signed("1101101101001110"),
    signed("0010010101100111"),
    signed("1101110100101000"),
    signed("0010000101111001"),
    signed("0010001001000110"),
    signed("0010010010111101"),
    signed("1101101010111110"),
    signed("1110001001000110"),
    signed("1110010000010001"),
    signed("0010010010111101"),
    signed("0001110000011111"),
    signed("1101101101101000"),
    signed("0001101101010000"));



constant lut_gs2i_data_58 : vector_of_signed16(0 to 63) := 
   (signed("1110000010010110"),
    signed("0010000111010110"),
    signed("0010001010001101"),
    signed("0010011110000010"),
    signed("1110100001110110"),
    signed("1101011111110011"),
    signed("1101001111001001"),
    signed("0010001110101110"),
    signed("0001100111110010"),
    signed("0010000010000001"),
    signed("1110001010101101"),
    signed("0010101101111001"),
    signed("0001110110010011"),
    signed("0001110100101110"),
    signed("0010001000100011"),
    signed("1110010101101000"),
    signed("1101001110101011"),
    signed("1101101100010111"),
    signed("0010100010011011"),
    signed("1101011111110011"),
    signed("0001100110101001"),
    signed("0010001000101011"),
    signed("1110011111111101"),
    signed("0010101011000001"),
    signed("1110000011101100"),
    signed("0001110010101110"),
    signed("0001011110101101"),
    signed("1110101110001011"),
    signed("1110100100001001"),
    signed("1101110100111001"),
    signed("1110010010001100"),
    signed("1101111001100001"),
    signed("1101100010010110"),
    signed("0010000111110110"),
    signed("1101110110111011"),
    signed("0010001111000101"),
    signed("1101110000010011"),
    signed("0001100000111101"),
    signed("0001111000000100"),
    signed("0010110010111100"),
    signed("0001111001011110"),
    signed("1101011110001001"),
    signed("0010110010111100"),
    signed("0010001110111010"),
    signed("1101011100111001"),
    signed("1110001010001000"),
    signed("1110100110000010"),
    signed("0001011011001100"),
    signed("0001110111101100"),
    signed("0010100010001110"),
    signed("1110110011010000"),
    signed("1101101000010111"),
    signed("0001111000111011"),
    signed("1101001101111011"),
    signed("0001110111110011"),
    signed("0001100011110010"),
    signed("0001110100101110"),
    signed("1101011110111100"),
    signed("1101111000000101"),
    signed("1110100111000111"),
    signed("0001110100101110"),
    signed("0001110100010101"),
    signed("1101000101110011"),
    signed("0001111010001011"));



constant lut_gs2i_data_59 : vector_of_signed16(0 to 63) := 
   (signed("1110100001101100"),
    signed("0001111101001110"),
    signed("0010001111011110"),
    signed("0010101110010001"),
    signed("1111001011100011"),
    signed("1101000011011001"),
    signed("1100110101110100"),
    signed("0010101011100111"),
    signed("0001101011010111"),
    signed("0001010101001110"),
    signed("1110011100100110"),
    signed("0011001111101000"),
    signed("0010000001110100"),
    signed("0001001110111000"),
    signed("0001101101101011"),
    signed("1110010111111101"),
    signed("1100110111111011"),
    signed("1110010000001011"),
    signed("0010110011110001"),
    signed("1101000011011001"),
    signed("0001100101111100"),
    signed("0010010001100011"),
    signed("1111000110010101"),
    signed("0010110101101000"),
    signed("1110001001000011"),
    signed("0001010011000100"),
    signed("0000101110110000"),
    signed("1111010011001001"),
    signed("1111000110010101"),
    signed("1110000001111110"),
    signed("1110011111100000"),
    signed("1101101010111001"),
    signed("1110000011010111"),
    signed("0001100010000001"),
    signed("1110011000100010"),
    signed("0010010110111110"),
    signed("1110010111110001"),
    signed("0001001010110100"),
    signed("0001111011000100"),
    signed("0010110111101111"),
    signed("0010000001110111"),
    signed("1110000011010111"),
    signed("0010110111101111"),
    signed("0001111100000001"),
    signed("1101000100101110"),
    signed("1110101011101110"),
    signed("1111001011100011"),
    signed("0000111001111010"),
    signed("0001001001011011"),
    signed("0010101110010001"),
    signed("1111100000001010"),
    signed("1101111000100001"),
    signed("0001001110111000"),
    signed("1100110000011000"),
    signed("0001100000000100"),
    signed("0000111011110001"),
    signed("0001001110111000"),
    signed("1101011011010010"),
    signed("1101100011100101"),
    signed("1111000000111001"),
    signed("0001001110111000"),
    signed("0001111000111101"),
    signed("1100101000110001"),
    signed("0010001101100001"));



constant lut_gs2i_data_60 : vector_of_signed16(0 to 63) := 
   (signed("1111001100001000"),
    signed("0001110001111010"),
    signed("0010010010101111"),
    signed("0010110101000011"),
    signed("1111110110010010"),
    signed("1100101111101001"),
    signed("1100101001010011"),
    signed("0011000011010101"),
    signed("0001110100101100"),
    signed("0000011100111011"),
    signed("1110110111110001"),
    signed("0011100100111011"),
    signed("0010001111111100"),
    signed("0000100010010101"),
    signed("0001000100101010"),
    signed("1110010101010000"),
    signed("1100101101111011"),
    signed("1111000011110100"),
    signed("0010111011001000"),
    signed("1100101111101001"),
    signed("0001101011000100"),
    signed("0010010110000111"),
    signed("1111101110011000"),
    signed("0010110100011111"),
    signed("1110001100110110"),
    signed("0000101010010101"),
    signed("1111111101000000"),
    signed("1111110111000111"),
    signed("1111101001011100"),
    signed("1110011101011100"),
    signed("1110101000000110"),
    signed("1101011101010110"),
    signed("1110110110001010"),
    signed("0000101111100001"),
    signed("1111000111001100"),
    signed("0010011100000010"),
    signed("1111001110100000"),
    signed("0000110001110001"),
    signed("0001111111010100"),
    signed("0010101111001111"),
    signed("0010001100101110"),
    signed("1110111011000110"),
    signed("0010101111001111"),
    signed("0001011011000001"),
    signed("1100110110101001"),
    signed("1111010100000011"),
    signed("1111110001010110"),
    signed("0000010111111100"),
    signed("0000010100000111"),
    signed("0010110000001000"),
    signed("0000001011011010"),
    signed("1110011001011000"),
    signed("0000011101011010"),
    signed("1100100000000001"),
    signed("0000111110101000"),
    signed("0000010001010100"),
    signed("0000100010010101"),
    signed("1101100000011001"),
    signed("1101010000110100"),
    signed("1111011011001110"),
    signed("0000100010010101"),
    signed("0001111111101001"),
    signed("1100011010010000"),
    signed("0010100001110110"));



constant lut_gs2i_data_61 : vector_of_signed16(0 to 63) := 
   (signed("1111111100101101"),
    signed("0001100111100100"),
    signed("0010010011110110"),
    signed("0010110011001100"),
    signed("0000011111011101"),
    signed("1100100110011011"),
    signed("1100101001100011"),
    signed("0011010011000000"),
    signed("0010000001001000"),
    signed("1111100000100011"),
    signed("1111011010011010"),
    signed("0011101100001100"),
    signed("0010011101011101"),
    signed("1111110011010001"),
    signed("0000010010100111"),
    signed("1110001110101111"),
    signed("1100110000001000"),
    signed("0000000000000000"),
    signed("0010111001011100"),
    signed("1100100110011011"),
    signed("0001110100011001"),
    signed("0010010110110111"),
    signed("0000010101101111"),
    signed("0010101010010010"),
    signed("1110001110101111"),
    signed("1111111100111000"),
    signed("1111001101100101"),
    signed("0000011000110111"),
    signed("0000001100000001"),
    signed("1111000100101011"),
    signed("1110101011000011"),
    signed("1101010011011010"),
    signed("1111110011001010"),
    signed("1111110111000111"),
    signed("1111111100111000"),
    signed("0010011101011101"),
    signed("0000001100110110"),
    signed("0000010101101111"),
    signed("0010000011111000"),
    signed("0010011101011101"),
    signed("0010010111101011"),
    signed("1111111100111000"),
    signed("0010011101011101"),
    signed("0000101111010011"),
    signed("1100110011010000"),
    signed("0000000000000000"),
    signed("0000010101101111"),
    signed("1111110110010010"),
    signed("1111011101100010"),
    signed("0010101001011110"),
    signed("0000110010011011"),
    signed("1111000110111111"),
    signed("1111101001100100"),
    signed("1100011101100001"),
    signed("0000010110011100"),
    signed("1111100111001001"),
    signed("1111110011010001"),
    signed("1101101011011101"),
    signed("1101000011000111"),
    signed("1111110110010010"),
    signed("1111110011010001"),
    signed("0010000111000000"),
    signed("1100011010011001"),
    signed("0010110011001100"));



constant lut_gs2i_data_62 : vector_of_signed16(0 to 63) := 
   (signed("0000101101110010"),
    signed("0001100000011000"),
    signed("0010010010101111"),
    signed("0010101010010000"),
    signed("0001000100100011"),
    signed("1100101000111111"),
    signed("1100110101011010"),
    signed("0011010111110110"),
    signed("0010001101010101"),
    signed("1110101000010000"),
    signed("0000000010010000"),
    signed("0011100100111011"),
    signed("0010100110110101"),
    signed("1111000110010011"),
    signed("1111011101110101"),
    signed("1110000110001011"),
    signed("1100111100111111"),
    signed("0000111100001100"),
    signed("0010110000010101"),
    signed("1100101000111111"),
    signed("0001111111100101"),
    signed("0010010100011100"),
    signed("0000111010001011"),
    signed("0010011010101000"),
    signed("1110001110100110"),
    signed("1111001111100110"),
    signed("1110100100101010"),
    signed("0000110111100001"),
    signed("0000101100110101"),
    signed("1111110100000010"),
    signed("1110101000000110"),
    signed("1101001111100100"),
    signed("0000110001100000"),
    signed("1111000000010010"),
    signed("0000110010101111"),
    signed("0010011010101111"),
    signed("0001001001110110"),
    signed("1111110110110010"),
    signed("0010000111101111"),
    signed("0010000111100001"),
    signed("0010011111111011"),
    signed("0000111110110110"),
    signed("0010000111100001"),
    signed("1111111101001111"),
    signed("1100111010010101"),
    signed("0000101011111101"),
    signed("0000110111001101"),
    signed("1111010101110010"),
    signed("1110101011111111"),
    signed("0010011100111010"),
    signed("0001010010111011"),
    signed("1111111100000101"),
    signed("1110111000111101"),
    signed("1100101000011011"),
    signed("1111101011000001"),
    signed("1111000000000101"),
    signed("1111000110010011"),
    signed("1101111001000011"),
    signed("1100111101100111"),
    signed("0000010010100000"),
    signed("1111000110010011"),
    signed("0010001101011111"),
    signed("1100101000000111"),
    signed("0010111101011110"));



constant lut_gs2i_data_63 : vector_of_signed16(0 to 63) := 
   (signed("0001011001100111"),
    signed("0001011110010110"),
    signed("0010001111011110"),
    signed("0010011100011011"),
    signed("0001100011011011"),
    signed("1100110111111011"),
    signed("1101001010111111"),
    signed("0011001111101100"),
    signed("0010010101110100"),
    signed("1101111011110101"),
    signed("0000101100101010"),
    signed("0011001111101000"),
    signed("0010101000110101"),
    signed("1110011111111100"),
    signed("1110101100111001"),
    signed("1101111101100101"),
    signed("1101010010010011"),
    signed("0001101111110101"),
    signed("0010100001111011"),
    signed("1100110111111011"),
    signed("0010001010000001"),
    signed("0010001111101011"),
    signed("0001011001101110"),
    signed("0010001001011010"),
    signed("1110001100011111"),
    signed("1110100111011100"),
    signed("1110000110000101"),
    signed("0001010010011011"),
    signed("0001001010110100"),
    signed("0000100111001101"),
    signed("1110011111100000"),
    signed("1101010011110101"),
    signed("0001101000001111"),
    signed("1110010010010101"),
    signed("0001100001111110"),
    signed("0010010011101010"),
    signed("0001111100101001"),
    signed("1111010101001111"),
    signed("0010001001111110"),
    signed("0001110010111010"),
    signed("0010100010100111"),
    signed("0001110111001001"),
    signed("0001110010111010"),
    signed("1111001001101001"),
    signed("1101001010111111"),
    signed("0001010100010010"),
    signed("0001010100100001"),
    signed("1110110111001100"),
    signed("1110000101010100"),
    signed("0010001101100001"),
    signed("0001101011000001"),
    signed("0000110010111011"),
    signed("1110010001000010"),
    signed("1100111111010010"),
    signed("1111000000000011"),
    signed("1110011110101011"),
    signed("1110011111111100"),
    signed("1110000101101111"),
    signed("1101000010110101"),
    signed("0000110000001101"),
    signed("1110011111111100"),
    signed("0010010001100100"),
    signed("1101000001011000"),
    signed("0010111101001011"));



constant lut_gs2i_data_64 : vector_of_signed16(0 to 63) := 
   (signed("0001111011000110"),
    signed("0001100010101101"),
    signed("0010001010001101"),
    signed("0010001100000111"),
    signed("0001111010100100"),
    signed("1101010010111000"),
    signed("1101100111111100"),
    signed("0010111001011101"),
    signed("0010010111100000"),
    signed("1101100001100101"),
    signed("0001010110110010"),
    signed("0010101101111001"),
    signed("0010100001000000"),
    signed("1110000100000000"),
    signed("1110000101111010"),
    signed("1101110110110000"),
    signed("1101101101100011"),
    signed("0010010011101001"),
    signed("0010010000100001"),
    signed("1101010010111000"),
    signed("0010010001011000"),
    signed("0010001001011101"),
    signed("0001110010111010"),
    signed("0001111010001111"),
    signed("1110001000101101"),
    signed("1110001000111000"),
    signed("1101110100110100"),
    signed("0001101001000101"),
    signed("0001100101001010"),
    signed("0001011001110000"),
    signed("1110010010001100"),
    signed("1101100001100000"),
    signed("0010001111101101"),
    signed("1101110011010001"),
    signed("0010000100101011"),
    signed("0010001000001101"),
    signed("0010011101101010"),
    signed("1110110001111001"),
    signed("0010001010000000"),
    signed("0001100100010110"),
    signed("0010011101010101"),
    signed("0010011101011101"),
    signed("0001100100010110"),
    signed("1110011001001011"),
    signed("1101100011101111"),
    signed("0001110101111000"),
    signed("0001101100110100"),
    signed("1110011011010000"),
    signed("1101101110001100"),
    signed("0001111110010111"),
    signed("0001111001001111"),
    signed("0001100110000001"),
    signed("1101110110010000"),
    signed("1101011111110111"),
    signed("1110011001000010"),
    signed("1110000100111110"),
    signed("1110000100000000"),
    signed("1110001110101010"),
    signed("1101010100001110"),
    signed("0001001111010101"),
    signed("1110000100000000"),
    signed("0010010010001000"),
    signed("1101100011100110"),
    signed("0010101111111110"));



-----------------------------------------------------------------
-----------------------------------------------------------------

GS2 q LUTs

constant lut_gs2q_data_1 : vector_of_signed16(0 to 63) := 
   (signed("1111111101110101"),
    signed("0010001100001001"),
    signed("0001101011100100"),
    signed("0010000001001010"),
    signed("0001111001100100"),
    signed("0010000111000001"),
    signed("1101111010101011"),
    signed("1110001011111010"),
    signed("0010010111101100"),
    signed("0010010010011000"),
    signed("1101011011010000"),
    signed("0001111011101011"),
    signed("0010000100010111"),
    signed("0010001011111100"),
    signed("1101110011000111"),
    signed("1101101011100010"),
    signed("1101110101001100"),
    signed("1110001110100100"),
    signed("0010100000011010"),
    signed("0001111100001110"),
    signed("1101111010101011"),
    signed("0010010110001010"),
    signed("0010000000100101"),
    signed("0010000010101011"),
    signed("0001101101101001"),
    signed("1110000101110111"),
    signed("1101111001100010"),
    signed("1101110000011101"),
    signed("0001111001000001"),
    signed("0001111101010111"),
    signed("0010000101010101"),
    signed("1110000011110010"),
    signed("1101111011000100"),
    signed("0010100100110000"),
    signed("1101100100111010"),
    signed("0010010100011110"),
    signed("0001111010101101"),
    signed("0010100101101110"),
    signed("1110001011111010"),
    signed("0010000101100000"),
    signed("0001100001010100"),
    signed("0010010000101100"),
    signed("0010101010000100"),
    signed("0001100001010100"),
    signed("1101110001111110"),
    signed("1110000100111010"),
    signed("0010001100010101"),
    signed("0010000001101101"),
    signed("1110000000100100"),
    signed("1101100111001011"),
    signed("0001101111111010"),
    signed("0001111110111001"),
    signed("0010001110100111"),
    signed("1101101101110011"),
    signed("1110001001101001"),
    signed("1101111011000100"),
    signed("1101110001111110"),
    signed("1101110011000111"),
    signed("1110010100000011"),
    signed("1101101111101101"),
    signed("0001101101000101"),
    signed("1101110011000111"),
    signed("0010010000110110"),
    signed("1110001001101001"));

constant lut_gs2q_data_2 : vector_of_signed16(0 to 63) := 
   (signed("1111111110001001"),
    signed("0010001111001100"),
    signed("0001111110100100"),
    signed("0001111011100000"),
    signed("0001101001100111"),
    signed("0010001011101001"),
    signed("1110100110010000"),
    signed("1110110001111001"),
    signed("0001101001110011"),
    signed("0001111110110000"),
    signed("1101110000010011"),
    signed("0010011111011000"),
    signed("0001001111101110"),
    signed("0001101100100110"),
    signed("1101110101010010"),
    signed("1101100011011010"),
    signed("1101110010110101"),
    signed("1110110000101011"),
    signed("0010010110110000"),
    signed("0001101101110100"),
    signed("1110100110010000"),
    signed("0010010101000110"),
    signed("0001111000100110"),
    signed("0010001111100101"),
    signed("0001100111110010"),
    signed("1101111101111011"),
    signed("1101110100111001"),
    signed("1101111011111000"),
    signed("0010001000101011"),
    signed("0010010000010110"),
    signed("0010101101001000"),
    signed("1101101111011111"),
    signed("1110011001000010"),
    signed("0010011110011011"),
    signed("1101101111010101"),
    signed("0010010010000001"),
    signed("0001100100101100"),
    signed("0010011001101110"),
    signed("1101100111111100"),
    signed("0001111111011011"),
    signed("0001100100010110"),
    signed("0001111001100110"),
    signed("0010011101101010"),
    signed("0001100100010110"),
    signed("1101010100010011"),
    signed("1110101001110001"),
    signed("0010011101010101"),
    signed("0010001100011010"),
    signed("1101101110100001"),
    signed("1101110111011001"),
    signed("0001100110101001"),
    signed("0001111001000010"),
    signed("0010110000001011"),
    signed("1101110110000011"),
    signed("1110110110111110"),
    signed("1101100001100000"),
    signed("1101101000100000"),
    signed("1101110101010010"),
    signed("1110001110101010"),
    signed("1110011010011101"),
    signed("0010001110101110"),
    signed("1101110101010010"),
    signed("0010000111010110"),
    signed("1110110011010000"));

constant lut_gs2q_data_3 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("0010000001110101"),
    signed("0010010011000001"),
    signed("0001110011100001"),
    signed("0001100000100000"),
    signed("0010001100000111"),
    signed("1111011000110011"),
    signed("1111010101001111"),
    signed("0000110000111010"),
    signed("0001100011011011"),
    signed("1110010111110001"),
    signed("0010111001001011"),
    signed("0000011010011010"),
    signed("0001000111010001"),
    signed("1110000011111111"),
    signed("1101110000111110"),
    signed("1101110101111111"),
    signed("1111001111110011"),
    signed("0001111010011111"),
    signed("0001100000100000"),
    signed("1111011000110011"),
    signed("0010001100001000"),
    signed("0001110100110110"),
    signed("0010010011101101"),
    signed("0001101011010111"),
    signed("1101111000001001"),
    signed("1110000001111110"),
    signed("1110011000010101"),
    signed("0010010001100011"),
    signed("0010011011010000"),
    signed("0011001000000101"),
    signed("1101011110000101"),
    signed("1111000000000011"),
    signed("0010000100001011"),
    signed("1110001010101111"),
    signed("0010000000001100"),
    signed("0001001100111011"),
    signed("0001110101000010"),
    signed("1101001010111111"),
    signed("0001111011000111"),
    signed("0001110010111010"),
    signed("0001010110011000"),
    signed("0001111100101001"),
    signed("0001110010111010"),
    signed("1100111111001110"),
    signed("1111001101101001"),
    signed("0010100010100111"),
    signed("0010010011101010"),
    signed("1101011111010101"),
    signed("1110010110011100"),
    signed("0001100101111100"),
    signed("0001100101100001"),
    signed("0011000010101011"),
    signed("1110001011100010"),
    signed("1111100010010000"),
    signed("1101010011110101"),
    signed("1101101010001100"),
    signed("1110000011111111"),
    signed("1110000101101111"),
    signed("1111001010111111"),
    signed("0010101011100111"),
    signed("1110000011111111"),
    signed("0001111101001110"),
    signed("1111100000001010"));

constant lut_gs2q_data_4 : vector_of_signed16(0 to 63) := 
   (signed("0000000000001010"),
    signed("0001100101011100"),
    signed("0010100111111011"),
    signed("0001101100011111"),
    signed("0001011100110110"),
    signed("0010000111111001"),
    signed("0000001011111110"),
    signed("1111110110110010"),
    signed("1111110100100010"),
    signed("0000111111100111"),
    signed("1111001110100000"),
    signed("0011001001101011"),
    signed("1111100110011000"),
    signed("0000011100100101"),
    signed("1110100000000011"),
    signed("1110010000011010"),
    signed("1101111011011111"),
    signed("1111101101100000"),
    signed("0001001101011000"),
    signed("0001010111111010"),
    signed("0000001011111110"),
    signed("0001111111010001"),
    signed("0001110011011111"),
    signed("0010010010100101"),
    signed("0001110100101100"),
    signed("1101110011000001"),
    signed("1110011101011100"),
    signed("1111000000100011"),
    signed("0010010110000111"),
    signed("0010100000011111"),
    signed("0011010111000001"),
    signed("1101001111101011"),
    signed("1111101011000001"),
    signed("0001010111110000"),
    signed("1110110101100110"),
    signed("0001011111000010"),
    signed("0000110001011100"),
    signed("0000111111001010"),
    signed("1100110101011010"),
    signed("0001110111001011"),
    signed("0010000111100001"),
    signed("0000101011101000"),
    signed("0001001001110110"),
    signed("0010000111100001"),
    signed("1100110101100000"),
    signed("1111110001000010"),
    signed("0010011111111011"),
    signed("0010010101110011"),
    signed("1101010101111010"),
    signed("1111000010100101"),
    signed("0001101011000100"),
    signed("0001000111111011"),
    signed("0011001000011110"),
    signed("1110101101111101"),
    signed("0000001011000110"),
    signed("1101001111100100"),
    signed("1101110010101011"),
    signed("1110100000000011"),
    signed("1101111001000011"),
    signed("1111111111010100"),
    signed("0011000011010101"),
    signed("1110100000000011"),
    signed("0001110001111010"),
    signed("0000001011011010"));

constant lut_gs2q_data_5 : vector_of_signed16(0 to 63) := 
   (signed("0000000001100100"),
    signed("0000111100111001"),
    signed("0010111001011100"),
    signed("0001100111100100"),
    signed("0001011110101010"),
    signed("0010000001001000"),
    signed("0000111011010101"),
    signed("0000010101101111"),
    signed("1110111010111110"),
    signed("0000010101101111"),
    signed("0000001100110110"),
    signed("0011001111111000"),
    signed("1110110111110110"),
    signed("1111110000001001"),
    signed("1111000110111111"),
    signed("1110111110000110"),
    signed("1110000001111001"),
    signed("0000001001101110"),
    signed("0000010101101111"),
    signed("0001010100111101"),
    signed("0000111011010101"),
    signed("0001110001010001"),
    signed("0001110100011001"),
    signed("0010001101111110"),
    signed("0010000001001000"),
    signed("1101101111010010"),
    signed("1111000100101011"),
    signed("1111110000001001"),
    signed("0010010110110111"),
    signed("0010100000100101"),
    signed("0011011001100101"),
    signed("1101000110100100"),
    signed("0000010110011100"),
    signed("0000011111011101"),
    signed("1111101010010001"),
    signed("0000110010011011"),
    signed("0000010010100111"),
    signed("0000000000000000"),
    signed("1100101001100011"),
    signed("0001110100011001"),
    signed("0010011101011101"),
    signed("1111111100111000"),
    signed("0000001100110110"),
    signed("0010011101011101"),
    signed("1100110110101110"),
    signed("0000010010100111"),
    signed("0010010111101011"),
    signed("0010010011101111"),
    signed("1101010010101101"),
    signed("1111110110010010"),
    signed("0001110100011001"),
    signed("0000100010011110"),
    signed("0011000011001001"),
    signed("1111011001100110"),
    signed("0000101111010011"),
    signed("1101010011011010"),
    signed("1101111110111000"),
    signed("1111000110111111"),
    signed("1101101011011101"),
    signed("0000110010011011"),
    signed("0011010011000000"),
    signed("1111000110111111"),
    signed("0001100111100100"),
    signed("0000110010011011"));

constant lut_gs2q_data_6 : vector_of_signed16(0 to 63) := 
   (signed("0000000010111000"),
    signed("0000001100001000"),
    signed("0011000011100010"),
    signed("0001100101110100"),
    signed("0001100101010000"),
    signed("0001111010001000"),
    signed("0001100010100100"),
    signed("0000110001110001"),
    signed("1110001010101010"),
    signed("1111101000111100"),
    signed("0001001001110110"),
    signed("0011001011011011"),
    signed("1110010010110000"),
    signed("1111000101111111"),
    signed("1111110101011011"),
    signed("1111110100110111"),
    signed("1110000111100110"),
    signed("0000100100110010"),
    signed("1111011011001010"),
    signed("0001010111111010"),
    signed("0001100010100100"),
    signed("0001100101010100"),
    signed("0001110111001011"),
    signed("0010000111110010"),
    signed("0010001101010101"),
    signed("1101101101100101"),
    signed("1111110100000010"),
    signed("0000100010000001"),
    signed("0010010100011100"),
    signed("0010011100010110"),
    signed("0011010000010111"),
    signed("1101000100111000"),
    signed("0000111110101000"),
    signed("1111100011000101"),
    signed("0000100001110111"),
    signed("1111111111010100"),
    signed("1111110001000010"),
    signed("1111000000110110"),
    signed("1100101001010011"),
    signed("0001110011011111"),
    signed("0010101111001111"),
    signed("1111001110010011"),
    signed("1111001110100000"),
    signed("0010101111001111"),
    signed("1101000001100111"),
    signed("0000110001011100"),
    signed("0010001100101110"),
    signed("0010001110101100"),
    signed("1101010101111010"),
    signed("0000101011001010"),
    signed("0001111111100101"),
    signed("1111110111111111"),
    signed("0010110101010001"),
    signed("0000001001111111"),
    signed("0001001101001011"),
    signed("1101011101010110"),
    signed("1110001011010100"),
    signed("1111110101011011"),
    signed("1101100000011001"),
    signed("0001011111000010"),
    signed("0011010111110110"),
    signed("1111110101011011"),
    signed("0001100000011000"),
    signed("0001010010111011"));

constant lut_gs2q_data_7 : vector_of_signed16(0 to 63) := 
   (signed("0000000011110011"),
    signed("1111010111101111"),
    signed("0011000010101011"),
    signed("0001101000000011"),
    signed("0001101111011010"),
    signed("0001110101000011"),
    signed("0001111110000010"),
    signed("0001001010110100"),
    signed("1101101001010111"),
    signed("1110111100101001"),
    signed("0001111100101001"),
    signed("0010111100100111"),
    signed("1101111010011000"),
    signed("1110100010000010"),
    signed("0000100111011101"),
    signed("0000101110110100"),
    signed("1110001011001010"),
    signed("0000111111000111"),
    signed("1110100101100101"),
    signed("0001100000100000"),
    signed("0001111110000010"),
    signed("0001011110010110"),
    signed("0001111011000111"),
    signed("0010000001110111"),
    signed("0010010101110100"),
    signed("1101101110011100"),
    signed("0000100111001101"),
    signed("0001010000111110"),
    signed("0010001111101011"),
    signed("0010010100111000"),
    signed("0010111100100111"),
    signed("1101001100001111"),
    signed("0001100000000100"),
    signed("1110101010110010"),
    signed("0001010101001110"),
    signed("1111001010111111"),
    signed("1111001101101001"),
    signed("1110001010111110"),
    signed("1100110101110100"),
    signed("0001110100110110"),
    signed("0010110111101111"),
    signed("1110100100001000"),
    signed("1110010111110001"),
    signed("0010110111101111"),
    signed("1101010100011001"),
    signed("0001001100111011"),
    signed("0010000001110111"),
    signed("0010001000000100"),
    signed("1101011111010101"),
    signed("0001011010101010"),
    signed("0010001010000001"),
    signed("1111001011110000"),
    signed("0010100001111011"),
    signed("0000111010011110"),
    signed("0001100011011010"),
    signed("1101101010111001"),
    signed("1110010100101001"),
    signed("0000100111011101"),
    signed("1101011011010010"),
    signed("0010000000001100"),
    signed("0011001111101100"),
    signed("0000100111011101"),
    signed("0001011110010110"),
    signed("0001101011000001"));

constant lut_gs2q_data_8 : vector_of_signed16(0 to 63) := 
   (signed("0000000100000100"),
    signed("1110100100011001"),
    signed("0010110100011000"),
    signed("0001101110100100"),
    signed("0001111011100100"),
    signed("0001110011101001"),
    signed("0010001011000111"),
    signed("0001100000111101"),
    signed("1101011011010010"),
    signed("1110010100000110"),
    signed("0010011101101010"),
    signed("0010100100011001"),
    signed("1101110000111101"),
    signed("1110000111101111"),
    signed("0001011001000101"),
    signed("0001100110000101"),
    signed("1110001011100111"),
    signed("0001011000111001"),
    signed("1101111100000110"),
    signed("0001101101110100"),
    signed("0010001011000111"),
    signed("0001011110100001"),
    signed("0001111111011011"),
    signed("0001111101101011"),
    signed("0010010111100000"),
    signed("1101110010000100"),
    signed("0001011001110000"),
    signed("0001111000011101"),
    signed("0010001001011101"),
    signed("0010001011010111"),
    signed("0010100000001101"),
    signed("1101011101100101"),
    signed("0001110111110011"),
    signed("1101111101111111"),
    signed("0001111101110101"),
    signed("1110011010011101"),
    signed("1110101001110001"),
    signed("1101100110010010"),
    signed("1101001111001001"),
    signed("0001111000100110"),
    signed("0010110010111100"),
    signed("1110000010000000"),
    signed("1101110000010011"),
    signed("0010110010111100"),
    signed("1101101101000101"),
    signed("0001100100101100"),
    signed("0001111001011110"),
    signed("0010000001010101"),
    signed("1101101110100001"),
    signed("0001111111000011"),
    signed("0010010001011000"),
    signed("1110100001000110"),
    signed("0010001100010100"),
    signed("0001100110110001"),
    signed("0001110001000111"),
    signed("1101111001100001"),
    signed("1110011000001110"),
    signed("0001011001000101"),
    signed("1101011110111100"),
    signed("0010010010000001"),
    signed("0010111001011101"),
    signed("0001011001000101"),
    signed("0001100010101101"),
    signed("0001111001001111"));

constant lut_gs2q_data_9 : vector_of_signed16(0 to 63) := 
   (signed("0000000001010101"),
    signed("1101110100001010"),
    signed("0010010101100111"),
    signed("0001111011010000"),
    signed("0010001010001111"),
    signed("0001110100101001"),
    signed("0010000110011110"),
    signed("0001110110010111"),
    signed("1101100000001011"),
    signed("1101110100001111"),
    signed("0010100101101110"),
    signed("0010000110011100"),
    signed("1101110101001100"),
    signed("1101110111011101"),
    signed("0010001000101110"),
    signed("0010010111101100"),
    signed("1110000110011100"),
    signed("0001101111101111"),
    signed("1101100110001101"),
    signed("0001111100001110"),
    signed("0010000110011110"),
    signed("0001101000111010"),
    signed("0010000101100000"),
    signed("0001111110010011"),
    signed("0010010010011000"),
    signed("1101111010100000"),
    signed("0010000101010101"),
    signed("0010010111010011"),
    signed("0010000100111011"),
    signed("0001111110111000"),
    signed("0001111111011100"),
    signed("1101111011000100"),
    signed("0010000001100011"),
    signed("1101100100100001"),
    signed("0010010100011110"),
    signed("1101101111101101"),
    signed("1110000100111010"),
    signed("1101010101111100"),
    signed("1101110001111110"),
    signed("0010000000100101"),
    signed("0010011100100111"),
    signed("1101101000010100"),
    signed("1101011111100110"),
    signed("0010100000111101"),
    signed("1110000111100100"),
    signed("0001111010101101"),
    signed("0001110111010011"),
    signed("0001111001100100"),
    signed("1110000000100100"),
    signed("0010010110001011"),
    signed("0010010110001010"),
    signed("1101111000111111"),
    signed("0001110101001110"),
    signed("0010001001010010"),
    signed("0001110111111000"),
    signed("1110000100110000"),
    signed("1110010010010111"),
    signed("0010000100010111"),
    signed("1101101111010100"),
    signed("0010010100011110"),
    signed("0010010011010110"),
    signed("0010000100010111"),
    signed("0001101011100100"),
    signed("0001111010100011"));

constant lut_gs2q_data_10 : vector_of_signed16(0 to 63) := 
   (signed("0000000000001111"),
    signed("1101001111001001"),
    signed("0001101110001001"),
    signed("0010000110011111"),
    signed("0010010111001101"),
    signed("0001111010101101"),
    signed("0001110111001000"),
    signed("0010001000001101"),
    signed("1101111101111111"),
    signed("1101011100010111"),
    signed("0010011001101110"),
    signed("0001011110001010"),
    signed("1110001001000101"),
    signed("1101110101010010"),
    signed("0010101100011101"),
    signed("0010111101001011"),
    signed("1101111110101011"),
    signed("0010001001100100"),
    signed("1101100000001111"),
    signed("0010010000100001"),
    signed("0001110111001000"),
    signed("0001111010001011"),
    signed("0010001010000000"),
    signed("0010000001011001"),
    signed("0001111110110000"),
    signed("1110000100100000"),
    signed("0010101101001000"),
    signed("0010100101001100"),
    signed("0001111100010100"),
    signed("0001110111010111"),
    signed("0001010110000010"),
    signed("1110011100111101"),
    signed("0001111110110111"),
    signed("1101011111000000"),
    signed("0010011000110111"),
    signed("1101010100001110"),
    signed("1101100011101111"),
    signed("1101011110100111"),
    signed("1110100010100010"),
    signed("0010001001011101"),
    signed("0001110111101100"),
    signed("1101011010110000"),
    signed("1101100101010100"),
    signed("0001111011011011"),
    signed("1110100100110100"),
    signed("0010001000001101"),
    signed("0001111001010001"),
    signed("0001110100011001"),
    signed("1110011011010000"),
    signed("0010010110111110"),
    signed("0010010101000110"),
    signed("1101011000101101"),
    signed("0001100101101011"),
    signed("0010100010011011"),
    signed("0001110100110101"),
    signed("1110010001011100"),
    signed("1110000101110001"),
    signed("0010101000101111"),
    signed("1110001010001000"),
    signed("0010000100101011"),
    signed("0001100110000101"),
    signed("0010101000101111"),
    signed("0001111110100100"),
    signed("0001110101010011"));

constant lut_gs2q_data_11 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("1100110101110100"),
    signed("0000111010100001"),
    signed("0010010101000111"),
    signed("0010011110100101"),
    signed("0010000111010011"),
    signed("0001011000100100"),
    signed("0010010011101010"),
    signed("1110101010110010"),
    signed("1101001010111100"),
    signed("0001110101000010"),
    signed("0000110100011101"),
    signed("1110101100111100"),
    signed("1110000011111111"),
    signed("0011001000010101"),
    signed("0011010001110010"),
    signed("1101110111111100"),
    signed("0010011110100100"),
    signed("1101110000111010"),
    signed("0010100001111011"),
    signed("0001011000100100"),
    signed("0010001101100001"),
    signed("0010001001111110"),
    signed("0010000011111101"),
    signed("0001100011011011"),
    signed("1110001100011111"),
    signed("0011001000000101"),
    signed("0010101000110101"),
    signed("0001110110111101"),
    signed("0001101111011010"),
    signed("0000101100110111"),
    signed("1111000111101001"),
    signed("0001110010010100"),
    signed("1101101011011110"),
    signed("0010001100111100"),
    signed("1101000010110101"),
    signed("1101001010111111"),
    signed("1110000001010001"),
    signed("1111010110101100"),
    signed("0010001111101011"),
    signed("0001001001011011"),
    signed("1101011011010010"),
    signed("1101111101111011"),
    signed("0001001011100010"),
    signed("1111000110000110"),
    signed("0010010011101010"),
    signed("0001111100010111"),
    signed("0001110100110110"),
    signed("1110110111001100"),
    signed("0010000111101111"),
    signed("0010001100001000"),
    signed("1101000100101110"),
    signed("0001011000111001"),
    signed("0010110011110001"),
    signed("0001100101100001"),
    signed("1110010111111101"),
    signed("1101110110100110"),
    signed("0011000110001110"),
    signed("1110101011101110"),
    signed("0001100001111110"),
    signed("0000101110110100"),
    signed("0011000110001110"),
    signed("0010010011000001"),
    signed("0001100011011010"));

constant lut_gs2q_data_12 : vector_of_signed16(0 to 63) := 
   (signed("1111111101101100"),
    signed("1100101001010011"),
    signed("0000000001110101"),
    signed("0010100010101010"),
    signed("0010100001110010"),
    signed("0010010110000000"),
    signed("0000110000011010"),
    signed("0010011010101111"),
    signed("1111100011000101"),
    signed("1101000010011111"),
    signed("0000111111001010"),
    signed("0000001001101110"),
    signed("1111011010100111"),
    signed("1110100000000011"),
    signed("0011011000011001"),
    signed("0011010111100001"),
    signed("1101110001010100"),
    signed("0010101111010110"),
    signed("1110010011101000"),
    signed("0010110000010101"),
    signed("0000110000011010"),
    signed("0010100001110110"),
    signed("0010000111101111"),
    signed("0010000111011110"),
    signed("0000111111100111"),
    signed("1110010011100001"),
    signed("0011010111000001"),
    signed("0010100001111001"),
    signed("0001110011001010"),
    signed("0001101010001100"),
    signed("0000000011111110"),
    signed("1111110101101101"),
    signed("0001011010100001"),
    signed("1110001010010110"),
    signed("0001101111111010"),
    signed("1100111101100111"),
    signed("1100111010010101"),
    signed("1110110110011110"),
    signed("0000001100010010"),
    signed("0010010100011100"),
    signed("0000010100000111"),
    signed("1101100101010101"),
    signed("1110100111111100"),
    signed("0000010011110011"),
    signed("1111101000000100"),
    signed("0010011010101111"),
    signed("0010000001101101"),
    signed("0001111000011010"),
    signed("1111010101110010"),
    signed("0001101000000000"),
    signed("0001111111010001"),
    signed("1100111011100101"),
    signed("0001010010001010"),
    signed("0010111011001000"),
    signed("0001001100110111"),
    signed("1110011010001100"),
    signed("1101100101011000"),
    signed("0011011000101110"),
    signed("1111010100000011"),
    signed("0000110010101111"),
    signed("1111110100110111"),
    signed("0011011000101110"),
    signed("0010100111111011"),
    signed("0001001000001111"));

constant lut_gs2q_data_13 : vector_of_signed16(0 to 63) := 
   (signed("1111111100101101"),
    signed("1100101001100011"),
    signed("1111001010000111"),
    signed("0010101100100110"),
    signed("0010100000100101"),
    signed("0010100011101101"),
    signed("0000000011001000"),
    signed("0010011101011101"),
    signed("0000011111011101"),
    signed("1101000010101111"),
    signed("0000000000000000"),
    signed("1111100000100011"),
    signed("0000001100110110"),
    signed("1111000110111111"),
    signed("0011011011111001"),
    signed("0011001111111000"),
    signed("1101101100010001"),
    signed("0010111010001001"),
    signed("1111000011110111"),
    signed("0010111001011100"),
    signed("0000000011001000"),
    signed("0010110011001100"),
    signed("0010000011111000"),
    signed("0010001010110110"),
    signed("0000010101101111"),
    signed("1110011000011100"),
    signed("0011011001100101"),
    signed("0010010011101111"),
    signed("0001110001010001"),
    signed("0001101000011000"),
    signed("1111011101011011"),
    signed("0000100011010010"),
    signed("0000111001000001"),
    signed("1110110111110110"),
    signed("0001000101000010"),
    signed("1101000011000111"),
    signed("1100110011010000"),
    signed("1111110110010010"),
    signed("0000111110011101"),
    signed("0010010110110111"),
    signed("1111011101100010"),
    signed("1101110101001010"),
    signed("1111011101011011"),
    signed("1111011010011010"),
    signed("0000001001101110"),
    signed("0010011101011101"),
    signed("0010000111101110"),
    signed("0001111110000111"),
    signed("1111110110010010"),
    signed("0000111011010101"),
    signed("0001110001010001"),
    signed("1100111100111110"),
    signed("0001010001110101"),
    signed("0010111001011100"),
    signed("0000101100001011"),
    signed("1110011000011100"),
    signed("1101010101101110"),
    signed("0011011111000001"),
    signed("0000000000000000"),
    signed("1111111100111000"),
    signed("1110111110000110"),
    signed("0011011111000001"),
    signed("0010111001011100"),
    signed("0000100101100110"));

constant lut_gs2q_data_14 : vector_of_signed16(0 to 63) := 
   (signed("1111111100001101"),
    signed("1100110101011010"),
    signed("1110011001101101"),
    signed("0010110000011100"),
    signed("0010011011000011"),
    signed("0010101100111010"),
    signed("1111010101101011"),
    signed("0010011100000010"),
    signed("0001010111110000"),
    signed("1101001010111001"),
    signed("1111000000110110"),
    signed("1110111011011101"),
    signed("0000111101110000"),
    signed("1111110101011011"),
    signed("0011010010111110"),
    signed("0010111101100101"),
    signed("1101101010001101"),
    signed("0010111101001101"),
    signed("1111111011110001"),
    signed("0010111011001000"),
    signed("1111010101101011"),
    signed("0010111101011110"),
    signed("0001111111010100"),
    signed("0010001100110101"),
    signed("1111101000111100"),
    signed("1110011010001100"),
    signed("0011010000010111"),
    signed("0010000010100110"),
    signed("0001110001011010"),
    signed("0001101010001100"),
    signed("1110111011001001"),
    signed("0001001100010011"),
    signed("0000010000000001"),
    signed("1111101110110010"),
    signed("0000010000111001"),
    signed("1101010000110100"),
    signed("1100110110101001"),
    signed("0000110111010000"),
    signed("0001101000010100"),
    signed("0010010110000111"),
    signed("1110101011111111"),
    signed("1110000110011001"),
    signed("0000010111001011"),
    signed("1110100110001110"),
    signed("0000101010001110"),
    signed("0010011100000010"),
    signed("0010001100100000"),
    signed("0010000100100001"),
    signed("0000010111111100"),
    signed("0000000110100010"),
    signed("0001100101010100"),
    signed("1101000111101011"),
    signed("0001010111100110"),
    signed("0010110000010101"),
    signed("0000000101010101"),
    signed("1110010011100001"),
    signed("1101001011100001"),
    signed("0011011000101110"),
    signed("0000101011111101"),
    signed("1111000111001100"),
    signed("1110010000011010"),
    signed("0011011000101110"),
    signed("0011000011100010"),
    signed("1111111101110000"));

constant lut_gs2q_data_15 : vector_of_signed16(0 to 63) := 
   (signed("1111111100010110"),
    signed("1101001010111111"),
    signed("1101110110011010"),
    signed("0010101100001011"),
    signed("0010010001100011"),
    signed("0010101110010101"),
    signed("1110101100111100"),
    signed("0010010110111110"),
    signed("0010000100001011"),
    signed("1101011001110110"),
    signed("1110001010111110"),
    signed("1110011100100101"),
    signed("0001100111011110"),
    signed("0000100111011101"),
    signed("0010111110101000"),
    signed("0010100100000000"),
    signed("1101101100010110"),
    signed("0010110111001011"),
    signed("0000110101000001"),
    signed("0010110011110001"),
    signed("1110101100111100"),
    signed("0010111101001011"),
    signed("0001111011000100"),
    signed("0010001100000111"),
    signed("1110111100101001"),
    signed("1110010111111101"),
    signed("0010111100100111"),
    signed("0001110010111010"),
    signed("0001110011100001"),
    signed("0001101111011010"),
    signed("1110011110101011"),
    signed("0001101100111000"),
    signed("1111100010010000"),
    signed("0000101001010100"),
    signed("1111011000110011"),
    signed("1101100011100101"),
    signed("1101000100101110"),
    signed("0001101111110101"),
    signed("0010000101101000"),
    signed("0010010001100011"),
    signed("1110000101010100"),
    signed("1110010100101001"),
    signed("0001001101100111"),
    signed("1101111101101110"),
    signed("0001001000110100"),
    signed("0010010110111110"),
    signed("0010001110001101"),
    signed("0010001010000001"),
    signed("0000111001111010"),
    signed("1111001111000110"),
    signed("0001011110010110"),
    signed("1101011001111001"),
    signed("0001100010100110"),
    signed("0010100001111011"),
    signed("1111011010101010"),
    signed("1110001100011111"),
    signed("1101001010011000"),
    signed("0011000110001110"),
    signed("0001010100010010"),
    signed("1110011000100010"),
    signed("1101110000111110"),
    signed("0011000110001110"),
    signed("0011000010101011"),
    signed("1111010011010110"));

constant lut_gs2q_data_16 : vector_of_signed16(0 to 63) := 
   (signed("1111111101001100"),
    signed("1101100111111100"),
    signed("1101100100101000"),
    signed("0010011110100000"),
    signed("0010000100011111"),
    signed("0010100101011001"),
    signed("1110001101010010"),
    signed("0010001111000101"),
    signed("0010011110011011"),
    signed("1101101110010100"),
    signed("1101100110010010"),
    signed("1110000101011100"),
    signed("0010000100111000"),
    signed("0001011001000101"),
    signed("0010100000100111"),
    signed("0010000110100110"),
    signed("1101110011100110"),
    signed("0010100111010111"),
    signed("0001101001101111"),
    signed("0010100010011011"),
    signed("1110001101010010"),
    signed("0010101111111110"),
    signed("0001111000000100"),
    signed("0010000111011101"),
    signed("1110010100000110"),
    signed("1110010001011100"),
    signed("0010100000001101"),
    signed("0001101000100011"),
    signed("0001110111010011"),
    signed("0001110111010111"),
    signed("1110001001001011"),
    signed("0010000001110101"),
    signed("1110110010110010"),
    signed("0001100001101011"),
    signed("1110100010000100"),
    signed("1101111000000101"),
    signed("1101011100111001"),
    signed("0010010111110101"),
    signed("0010010011010000"),
    signed("0010001000101011"),
    signed("1101101110001100"),
    signed("1110011100011010"),
    signed("0001111001111001"),
    signed("1101100110000100"),
    signed("0001100100110000"),
    signed("0010001111000101"),
    signed("0010001011001011"),
    signed("0010001101001011"),
    signed("0001011011001100"),
    signed("1110011010011001"),
    signed("0001011110100001"),
    signed("1101110001011111"),
    signed("0001110001100010"),
    signed("0010010000100001"),
    signed("1110101110110110"),
    signed("1110000100100000"),
    signed("1101010100111111"),
    signed("0010101000101111"),
    signed("0001110101111000"),
    signed("1101110110111011"),
    signed("1101100011011010"),
    signed("0010101000101111"),
    signed("0010110100011000"),
    signed("1110101001001110"));

constant lut_gs2q_data_17 : vector_of_signed16(0 to 63) := 
   (signed("0000000000110110"),
    signed("1110000111100100"),
    signed("1101100100100001"),
    signed("0010000100111100"),
    signed("0001110110010111"),
    signed("0010010010111101"),
    signed("1101111100001100"),
    signed("0010000011001111"),
    signed("0010100000011010"),
    signed("1110000100111010"),
    signed("1101011010010010"),
    signed("1101110100101000"),
    signed("0010010000001000"),
    signed("0010000100010111"),
    signed("0001111001000001"),
    signed("0001101010011011"),
    signed("1110000010101001"),
    signed("0010010000000111"),
    signed("0010010010111101"),
    signed("0010001001010010"),
    signed("1101110111110110"),
    signed("0010010010111101"),
    signed("0001111001001011"),
    signed("0001111011101011"),
    signed("1101110100001111"),
    signed("1110000100110000"),
    signed("0001111011000110"),
    signed("0001101000010101"),
    signed("0001111110011111"),
    signed("0010000011001111"),
    signed("1101111101010101"),
    signed("0010001011001101"),
    signed("1110000110111111"),
    signed("0010010000101100"),
    signed("1101110011101011"),
    signed("1110001001000110"),
    signed("1101111111111111"),
    signed("0010100111011010"),
    signed("0010001101011110"),
    signed("0001111001000001"),
    signed("1101100111001011"),
    signed("1110011101101110"),
    signed("0010010100011110"),
    signed("1101100000001011"),
    signed("0001111111011100"),
    signed("0010000111100101"),
    signed("0010000100010111"),
    signed("0010001010110100"),
    signed("0001111000011100"),
    signed("1101101010111110"),
    signed("0001101000111010"),
    signed("1110001110100100"),
    signed("0010000000100101"),
    signed("0010000000100101"),
    signed("1110000010101001"),
    signed("1101111010100000"),
    signed("1101101010011001"),
    signed("0010000100010111"),
    signed("0010010000101100"),
    signed("1101101000110111"),
    signed("1101100111001011"),
    signed("0010000000000001"),
    signed("0010011001111101"),
    signed("1101111111111111"));

constant lut_gs2q_data_18 : vector_of_signed16(0 to 63) := 
   (signed("0000000010011110"),
    signed("1110101110001011"),
    signed("1101111100100100"),
    signed("0001100110111110"),
    signed("0001100100101100"),
    signed("0001110100100001"),
    signed("1101111001000101"),
    signed("0001110111010111"),
    signed("0010001011111110"),
    signed("1110011111001100"),
    signed("1101100010010110"),
    signed("1101110000101000"),
    signed("0010001110000101"),
    signed("0010101000101111"),
    signed("0001010001001010"),
    signed("0001001110110111"),
    signed("1110010110111011"),
    signed("0001101011111010"),
    signed("0010110000001011"),
    signed("0001100110110001"),
    signed("1101110101010110"),
    signed("0001101001111100"),
    signed("0001111000000100"),
    signed("0001101110101101"),
    signed("1101011100010111"),
    signed("1101111001100001"),
    signed("0001010010010011"),
    signed("0001101100011111"),
    signed("0010000101110100"),
    signed("0010001111000101"),
    signed("1101110100010111"),
    signed("0010000101100011"),
    signed("1101011011011110"),
    signed("0010110101010000"),
    signed("1101001010110000"),
    signed("1110011010110011"),
    signed("1110101001001110"),
    signed("0010011110111001"),
    signed("0001111011010101"),
    signed("0001101001000101"),
    signed("1101110111011001"),
    signed("1110010001101000"),
    signed("0010011100110011"),
    signed("1101110011001101"),
    signed("0010010001011111"),
    signed("0001111011000110"),
    signed("0001110010011100"),
    signed("0010001001010000"),
    signed("0010010010111011"),
    signed("1101001010111101"),
    signed("0001111010001011"),
    signed("1110101100101111"),
    signed("0010010000100001"),
    signed("0001110001100010"),
    signed("1101011011101011"),
    signed("1101110010000100"),
    signed("1110001100101101"),
    signed("0001011001000101"),
    signed("0010100001000100"),
    signed("1101101001110010"),
    signed("1110000010001011"),
    signed("0001010101010111"),
    signed("0001110001110111"),
    signed("1101011100111001"));

constant lut_gs2q_data_19 : vector_of_signed16(0 to 63) := 
   (signed("0000000011110001"),
    signed("1111010011001001"),
    signed("1110100011011111"),
    signed("0000111111111101"),
    signed("0001001100111011"),
    signed("0001001001011000"),
    signed("1110000001111110"),
    signed("0001101111011010"),
    signed("0001100110001000"),
    signed("1110111110110011"),
    signed("1110000011010111"),
    signed("1101110001110011"),
    signed("0001111000100101"),
    signed("0011000110001110"),
    signed("0000100101010110"),
    signed("0000110010010011"),
    signed("1110101101100101"),
    signed("0001000011010111"),
    signed("0011000010101011"),
    signed("0000111010011110"),
    signed("1101111111111000"),
    signed("0000111010100001"),
    signed("0001111011000100"),
    signed("0001011001101110"),
    signed("1101001010111100"),
    signed("1101101010111001"),
    signed("0000101010110001"),
    signed("0001111010100000"),
    signed("0010001001111110"),
    signed("0010010110111110"),
    signed("1101110011111001"),
    signed("0001101110111110"),
    signed("1100111001110010"),
    signed("0011001111101100"),
    signed("1100110000010100"),
    signed("1110100101000000"),
    signed("1111010011010110"),
    signed("0010000010000101"),
    signed("0001011000100100"),
    signed("0001010010011011"),
    signed("1110010110011100"),
    signed("1110000000010011"),
    signed("0010010100100010"),
    signed("1110010110011100"),
    signed("0010100000101011"),
    signed("0001110001100000"),
    signed("0001011011110101"),
    signed("0010000010011011"),
    signed("0010101011100111"),
    signed("1100110101110100"),
    signed("0010001101100001"),
    signed("1111001000001101"),
    signed("0010100001111011"),
    signed("0001100010100110"),
    signed("1100111111010010"),
    signed("1101101110011100"),
    signed("1110111100000101"),
    signed("0000100111011101"),
    signed("0010100100101110"),
    signed("1101111111110100"),
    signed("1110101010110010"),
    signed("0000100101010110"),
    signed("0000111100101000"),
    signed("1101000100101110"));

constant lut_gs2q_data_20 : vector_of_signed16(0 to 63) := 
   (signed("0000000100011111"),
    signed("1111110111000111"),
    signed("1111010110100011"),
    signed("0000010100111111"),
    signed("0000110001011100"),
    signed("0000010111010101"),
    signed("1110011000100000"),
    signed("0001101010001100"),
    signed("0000110001110100"),
    signed("1111100000011110"),
    signed("1110110110001010"),
    signed("1101111000011011"),
    signed("0001010100010110"),
    signed("0011011000101110"),
    signed("1111111010101011"),
    signed("0000010111001000"),
    signed("1111001000011111"),
    signed("0000010111000100"),
    signed("0011001000011110"),
    signed("0000001001111111"),
    signed("1110011000110101"),
    signed("0000000110110001"),
    signed("0001111111010100"),
    signed("0000111111000111"),
    signed("1101000010011111"),
    signed("1101011101010110"),
    signed("0000000100010010"),
    signed("0010001101010010"),
    signed("0010001100101010"),
    signed("0010011100000010"),
    signed("1101111000000111"),
    signed("0001001011111110"),
    signed("1100100010010110"),
    signed("0011011100110001"),
    signed("1100100011001111"),
    signed("1110101001001111"),
    signed("1111111101110000"),
    signed("0001010011001001"),
    signed("0000101011011110"),
    signed("0000110111100001"),
    signed("1111000010100101"),
    signed("1101101010110100"),
    signed("0001111010100110"),
    signed("1111000111100000"),
    signed("0010101010000110"),
    signed("0001101001111000"),
    signed("0000111110110010"),
    signed("0001111001110101"),
    signed("0010111110011001"),
    signed("1100101110001111"),
    signed("0010100001110110"),
    signed("1111100010110100"),
    signed("0010110000010101"),
    signed("0001010111100110"),
    signed("1100101101010111"),
    signed("1101101101100101"),
    signed("1111110001111110"),
    signed("1111110101011011"),
    signed("0010011111100111"),
    signed("1110100101111010"),
    signed("1111011110001001"),
    signed("1111110101101111"),
    signed("0000000001100001"),
    signed("1100110110101001"));

constant lut_gs2q_data_21 : vector_of_signed16(0 to 63) := 
   (signed("0000000100011101"),
    signed("0000011000110111"),
    signed("0000001111001001"),
    signed("1111101001100100"),
    signed("0000010010100111"),
    signed("1111100011010100"),
    signed("1110111010111110"),
    signed("0001101000011000"),
    signed("1111110110010010"),
    signed("0000000011001000"),
    signed("1111110011001010"),
    signed("1110000010000000"),
    signed("0000100101100110"),
    signed("0011011111000001"),
    signed("1111010011110101"),
    signed("1111111100111000"),
    signed("1111100111001001"),
    signed("1111101010010001"),
    signed("0011000011001001"),
    signed("1111011001100110"),
    signed("1110111110000110"),
    signed("1111010011110101"),
    signed("0010000011111000"),
    signed("0000011111011101"),
    signed("1101000010101111"),
    signed("1101010011011010"),
    signed("1111100000100011"),
    signed("0010100000100101"),
    signed("0010001101100110"),
    signed("0010011101011101"),
    signed("1101111110111000"),
    signed("0000100000001010"),
    signed("1100010111010001"),
    signed("0011011100101101"),
    signed("1100100011010011"),
    signed("1110100111100110"),
    signed("0000100101100110"),
    signed("0000011000110111"),
    signed("1111111001011010"),
    signed("0000011000110111"),
    signed("1111110110010010"),
    signed("1101010101101110"),
    signed("0001010001111000"),
    signed("0000000000000000"),
    signed("0010101101010011"),
    signed("0001100101010000"),
    signed("0000011100010101"),
    signed("0001110001010001"),
    signed("0011001001010010"),
    signed("1100110011010000"),
    signed("0010110011001100"),
    signed("1111111100111000"),
    signed("0010111001011100"),
    signed("0001010001110101"),
    signed("1100100111001111"),
    signed("1101101111010010"),
    signed("0000101000101110"),
    signed("1111000110111111"),
    signed("0010010100100011"),
    signed("1111010111010010"),
    signed("0000010101101111"),
    signed("1111001010000111"),
    signed("1111000110111111"),
    signed("1100110011010000"));

constant lut_gs2q_data_22 : vector_of_signed16(0 to 63) := 
   (signed("0000000011100111"),
    signed("0000110111100001"),
    signed("0001000101110011"),
    signed("1111000001011000"),
    signed("1111110001000010"),
    signed("1110110010111001"),
    signed("1111100110101100"),
    signed("0001101010001100"),
    signed("1110111011111010"),
    signed("0000100101100111"),
    signed("0000110001100000"),
    signed("1110001011101001"),
    signed("1111110001101001"),
    signed("0011011000101110"),
    signed("1110110011001001"),
    signed("1111100010110100"),
    signed("0000001000111001"),
    signed("1111000000011001"),
    signed("0010110101010001"),
    signed("1110101101111101"),
    signed("1111101100011100"),
    signed("1110100111000011"),
    signed("0010000111101111"),
    signed("1111111011101110"),
    signed("1101001010111001"),
    signed("1101001111100100"),
    signed("1111000000111001"),
    signed("0010101111100100"),
    signed("0010001100101010"),
    signed("0010011010101111"),
    signed("1110000101111000"),
    signed("1111101111111100"),
    signed("1100011001111100"),
    signed("0011010000101011"),
    signed("1100101111010101"),
    signed("1110100000110100"),
    signed("0001001000001111"),
    signed("1111011011011111"),
    signed("1111001000010101"),
    signed("1111110111000111"),
    signed("0000101011001010"),
    signed("1101000110000101"),
    signed("0000011110100100"),
    signed("0000111000100000"),
    signed("0010101010000110"),
    signed("0001100100011100"),
    signed("1111110101111110"),
    signed("0001101010110000"),
    signed("0011001010100000"),
    signed("1101000010110000"),
    signed("0010111101011110"),
    signed("0000010111001000"),
    signed("0010111011001000"),
    signed("0001010010001010"),
    signed("1100101101010111"),
    signed("1101110011000001"),
    signed("0001011010000110"),
    signed("1110100000000011"),
    signed("0010000110111101"),
    signed("0000001110000010"),
    signed("0001001010011010"),
    signed("1110100101110011"),
    signed("1110010011111101"),
    signed("1100111010010101"));

constant lut_gs2q_data_23 : vector_of_signed16(0 to 63) := 
   (signed("0000000010000011"),
    signed("0001010010011011"),
    signed("0001110011001011"),
    signed("1110011111111100"),
    signed("1111001101101001"),
    signed("1110001011100010"),
    signed("0000011000010011"),
    signed("0001101111011010"),
    signed("1110001010111110"),
    signed("0001000110101101"),
    signed("0001101000001111"),
    signed("1110010010100011"),
    signed("1110111110001011"),
    signed("0011000110001110"),
    signed("1110011010011111"),
    signed("1111001000001101"),
    signed("0000101100110111"),
    signed("1110011100100101"),
    signed("0010100001111011"),
    signed("1110001011100010"),
    signed("0000011111111010"),
    signed("1110000101010100"),
    signed("0010001001111110"),
    signed("1111010101001111"),
    signed("1101011001110110"),
    signed("1101010011110101"),
    signed("1110100110010010"),
    signed("0010110101101000"),
    signed("0010001001111110"),
    signed("0010010011101010"),
    signed("1110001010111101"),
    signed("1111000000000011"),
    signed("1100101010111000"),
    signed("0010111010100001"),
    signed("1101000101011111"),
    signed("1110010110000110"),
    signed("0001100011011010"),
    signed("1110100011011111"),
    signed("1110011110000010"),
    signed("1111010011001001"),
    signed("0001011010101010"),
    signed("1101000000101011"),
    signed("1111100101100110"),
    signed("0001101001100100"),
    signed("0010100000101011"),
    signed("0001100111110011"),
    signed("1111001101101001"),
    signed("0001101000000011"),
    signed("0011000000110010"),
    signed("1101011001111001"),
    signed("0010111101001011"),
    signed("0000110010010011"),
    signed("0010110011110001"),
    signed("0001011000111001"),
    signed("1100111111010010"),
    signed("1101111000001001"),
    signed("0010000000001100"),
    signed("1110000011111111"),
    signed("0001111010010001"),
    signed("0001000011111011"),
    signed("0001110101010001"),
    signed("1110001011100101"),
    signed("1101101110110100"),
    signed("1101001010111111"));

constant lut_gs2q_data_24 : vector_of_signed16(0 to 63) := 
   (signed("1111111111111110"),
    signed("0001101001000101"),
    signed("0010010001001001"),
    signed("1110001000001101"),
    signed("1110101001110001"),
    signed("1101110001110110"),
    signed("0001001100000000"),
    signed("0001110111010111"),
    signed("1101101010011110"),
    signed("0001100101001110"),
    signed("0010001111101101"),
    signed("1110010100011111"),
    signed("1110010000011100"),
    signed("0010101000101111"),
    signed("1110001011001011"),
    signed("1110101100101111"),
    signed("0001010001110101"),
    signed("1110000001010000"),
    signed("0010001100010100"),
    signed("1101110110000011"),
    signed("0001010100001000"),
    signed("1101110010011000"),
    signed("0010001010000000"),
    signed("1110101101101101"),
    signed("1101101110010100"),
    signed("1101100001100000"),
    signed("1110010001010011"),
    signed("0010101111001101"),
    signed("0010000101110100"),
    signed("0010001000001101"),
    signed("1110001100010111"),
    signed("1110010100110101"),
    signed("1101001001100001"),
    signed("0010011100011110"),
    signed("1101100011100010"),
    signed("1110001000110110"),
    signed("0001110101010011"),
    signed("1101111000010111"),
    signed("1101111111100010"),
    signed("1110101110001011"),
    signed("0001111111000011"),
    signed("1101001001001000"),
    signed("1110101100000101"),
    signed("0010001100110011"),
    signed("0010010001011111"),
    signed("0001101111001111"),
    signed("1110100101100100"),
    signed("0001101010011000"),
    signed("0010101011101101"),
    signed("1101110101101100"),
    signed("0010101111111110"),
    signed("0001001110110111"),
    signed("0010100010011011"),
    signed("0001100101101011"),
    signed("1101011011101011"),
    signed("1101111101111011"),
    signed("0010010110001110"),
    signed("1101110101010010"),
    signed("0001110001010110"),
    signed("0001110011010011"),
    signed("0010010000101011"),
    signed("1101111101011011"),
    signed("1101011100100000"),
    signed("1101100011101111"));

constant lut_gs2q_data_25 : vector_of_signed16(0 to 63) := 
   (signed("1111111011011101"),
    signed("0001111001000001"),
    signed("0010011001011010"),
    signed("1101111010000111"),
    signed("1110000100111010"),
    signed("1101101011001001"),
    signed("0010000000000001"),
    signed("0001111110111000"),
    signed("1101011100111100"),
    signed("0010000010000110"),
    signed("0010100000011010"),
    signed("1110001110000001"),
    signed("1101101010011001"),
    signed("0010000100010111"),
    signed("1110001000001000"),
    signed("1110010010111011"),
    signed("0001111000011100"),
    signed("1101101101101000"),
    signed("0001110101001110"),
    signed("1101110010001001"),
    signed("0010000010101011"),
    signed("1101101110001100"),
    signed("0010000101100000"),
    signed("1110000100111010"),
    signed("1110001001010000"),
    signed("1101111011000100"),
    signed("1110000100010101"),
    signed("0010011000010001"),
    signed("0001111110011111"),
    signed("0001110110010111"),
    signed("1110001011010111"),
    signed("1101110100000011"),
    signed("1101110001111110"),
    signed("0001111011000110"),
    signed("1110000100111010"),
    signed("1101111000011011"),
    signed("0001111010100011"),
    signed("1101100001110111"),
    signed("1101101110001100"),
    signed("1110000111100100"),
    signed("0010010001110100"),
    signed("1101011111000011"),
    signed("1101110100101000"),
    signed("0010011111110101"),
    signed("0001111111011100"),
    signed("0001110111111000"),
    signed("1101111101111010"),
    signed("0001110100010000"),
    signed("0010001110000010"),
    signed("1110010001001110"),
    signed("0010010010111101"),
    signed("0001101010011011"),
    signed("0010001001010010"),
    signed("0001111001100100"),
    signed("1110000010101001"),
    signed("1110000101110111"),
    signed("0010011011011111"),
    signed("1101110111011101"),
    signed("0001110000010011"),
    signed("0010010101100111"),
    signed("0010011011000110"),
    signed("1101111010000111"),
    signed("1101100001110111"),
    signed("1110000000100100"));

constant lut_gs2q_data_26 : vector_of_signed16(0 to 63) := 
   (signed("1111111001100000"),
    signed("0010001000101011"),
    signed("0010010001001001"),
    signed("1101111101011011"),
    signed("1101100011101111"),
    signed("1101110001110110"),
    signed("0010101101111001"),
    signed("0010001011010111"),
    signed("1101100110101111"),
    signed("0010011001100111"),
    signed("0010011010101100"),
    signed("1110000101110001"),
    signed("1101010001010000"),
    signed("0001011001000101"),
    signed("1110001110111001"),
    signed("1101110101001110"),
    signed("0010011000000100"),
    signed("1101101000100000"),
    signed("0001100101101011"),
    signed("1101111001111111"),
    signed("0010101110010111"),
    signed("1101111111100010"),
    signed("0001111111011011"),
    signed("1101011111110011"),
    signed("1110100010111011"),
    signed("1110011001000010"),
    signed("1101111000100011"),
    signed("0001110111101100"),
    signed("0001110111010011"),
    signed("0001100000111101"),
    signed("1110000101010011"),
    signed("1101011001011000"),
    signed("1110100011111101"),
    signed("0001010110000010"),
    signed("1110101001111110"),
    signed("1101101100111111"),
    signed("0001111001001111"),
    signed("1101100000001111"),
    signed("1101110010011000"),
    signed("1101100111111100"),
    signed("0010010011010000"),
    signed("1110001000100001"),
    signed("1101001001111111"),
    signed("0010011001111100"),
    signed("0001100100110000"),
    signed("0010000111001010"),
    signed("1101011011100111"),
    signed("0001111110010111"),
    signed("0001100110110101"),
    signed("1110110001001001"),
    signed("0001101001111100"),
    signed("0010000110100110"),
    signed("0001100110110001"),
    signed("0010010000000011"),
    signed("1110101110110110"),
    signed("1110001000101101"),
    signed("0010001100110011"),
    signed("1110000111101111"),
    signed("0001110101000100"),
    signed("0010101011000001"),
    signed("0010001100101111"),
    signed("1110001000001101"),
    signed("1101111100000110"),
    signed("1110100110000010"));

constant lut_gs2q_data_27 : vector_of_signed16(0 to 63) := 
   (signed("1111111000011100"),
    signed("0010010001100011"),
    signed("0001110011001011"),
    signed("1110001011100101"),
    signed("1101001010111111"),
    signed("1110001011100010"),
    signed("0011001111101000"),
    signed("0010010100111000"),
    signed("1110001000110111"),
    signed("0010101000010001"),
    signed("0010000010000101"),
    signed("1101110110100110"),
    signed("1101001000010001"),
    signed("0000100111011101"),
    signed("1110011100100110"),
    signed("1101011100000000"),
    signed("0010110101000001"),
    signed("1101101010001100"),
    signed("0001011000111001"),
    signed("1110010011001000"),
    signed("0011001101100010"),
    signed("1110011110000010"),
    signed("0001111011000111"),
    signed("1101000011011001"),
    signed("1111000000111001"),
    signed("1111000000000011"),
    signed("1101110011111001"),
    signed("0001001001011011"),
    signed("0001110011100001"),
    signed("0001001010110100"),
    signed("1101111000101101"),
    signed("1101001100001111"),
    signed("1111011110000000"),
    signed("0000101100110111"),
    signed("1111010011001001"),
    signed("1101100001011011"),
    signed("0001101011000001"),
    signed("1101110000111010"),
    signed("1110000101010100"),
    signed("1101001010111111"),
    signed("0010000101101000"),
    signed("1110111100000101"),
    signed("1100101000110001"),
    signed("0010000010010010"),
    signed("0001001000110100"),
    signed("0010010100111000"),
    signed("1101000011011001"),
    signed("0010001101100001"),
    signed("0000110110010111"),
    signed("1111001101101101"),
    signed("0000111010100001"),
    signed("0010100100000000"),
    signed("0000111010011110"),
    signed("0010100100000001"),
    signed("1111011010101010"),
    signed("1110001100011111"),
    signed("0001101001100100"),
    signed("1110100010000010"),
    signed("0001111100010111"),
    signed("0010110101101000"),
    signed("0001101101101011"),
    signed("1110011111111100"),
    signed("1110100101100101"),
    signed("1111001011100011"));

constant lut_gs2q_data_28 : vector_of_signed16(0 to 63) := 
   (signed("1111111000011110"),
    signed("0010010110000111"),
    signed("0001000101110011"),
    signed("1110100101110011"),
    signed("1100111010010101"),
    signed("1110110010111001"),
    signed("0011100100111011"),
    signed("0010011100010110"),
    signed("1110111100001111"),
    signed("0010101111110111"),
    signed("0001011000000100"),
    signed("1101100101011000"),
    signed("1101001011110101"),
    signed("1111110101011011"),
    signed("1110110010110101"),
    signed("1101000111010111"),
    signed("0011001010100110"),
    signed("1101110010101011"),
    signed("0001010010001010"),
    signed("1110111000101001"),
    signed("0011100000010100"),
    signed("1111001000010101"),
    signed("0001110111001011"),
    signed("1100101111101001"),
    signed("1111100000001010"),
    signed("1111101011000001"),
    signed("1101110011001011"),
    signed("0000010100000111"),
    signed("0001110001011010"),
    signed("0000110001110001"),
    signed("1101101010000000"),
    signed("1101001001110100"),
    signed("0000011000110100"),
    signed("0000000011111110"),
    signed("1111111100000010"),
    signed("1101011001010010"),
    signed("0001010010111011"),
    signed("1110010011101000"),
    signed("1110100111000011"),
    signed("1100110101011010"),
    signed("0001101000010100"),
    signed("1111110110111001"),
    signed("1100010101010101"),
    signed("0001011001110010"),
    signed("0000101010001110"),
    signed("0010100001010010"),
    signed("1100110100100101"),
    signed("0010011100111010"),
    signed("0000000010110001"),
    signed("1111101000111000"),
    signed("0000000110110001"),
    signed("0010111101100101"),
    signed("0000001001111111"),
    signed("0010110100111100"),
    signed("0000000101010101"),
    signed("1110001110100110"),
    signed("0000111000100000"),
    signed("1111000101111111"),
    signed("0010000110101001"),
    signed("0010110100011111"),
    signed("0000111111101110"),
    signed("1111000001011000"),
    signed("1111011011001010"),
    signed("1111110001010110"));

constant lut_gs2q_data_29 : vector_of_signed16(0 to 63) := 
   (signed("1111111001101001"),
    signed("0010010110110111"),
    signed("0000001111001001"),
    signed("1111001010000111"),
    signed("1100110011010000"),
    signed("1111100011010100"),
    signed("0011101100001100"),
    signed("0010100000100101"),
    signed("1111111001011010"),
    signed("0010110000011011"),
    signed("0000100010100101"),
    signed("1101010101101110"),
    signed("1101011000110110"),
    signed("1111000110111111"),
    signed("1111010000101101"),
    signed("1100111001110110"),
    signed("0011010110011101"),
    signed("1101111110111000"),
    signed("0001010001110101"),
    signed("1111100110011100"),
    signed("0011100101100111"),
    signed("1111111001011010"),
    signed("0001110100011001"),
    signed("1100100110011011"),
    signed("0000000000000000"),
    signed("0000010110011100"),
    signed("1101110101001010"),
    signed("1111011101100010"),
    signed("0001110001010001"),
    signed("0000010101101111"),
    signed("1101011100010011"),
    signed("1101010000010010"),
    signed("0001001110110000"),
    signed("1111011101011011"),
    signed("0000100010100101"),
    signed("1101010101101110"),
    signed("0000110010011011"),
    signed("1111000011110111"),
    signed("1111010011110101"),
    signed("1100101001100011"),
    signed("0000111110011101"),
    signed("0000110010011011"),
    signed("1100010000101100"),
    signed("0000100101100110"),
    signed("0000001001101110"),
    signed("0010101010010010"),
    signed("1100110000001000"),
    signed("0010101001011110"),
    signed("1111010000101101"),
    signed("0000000011001000"),
    signed("1111010011110101"),
    signed("0011001111111000"),
    signed("1111011001100110"),
    signed("0011000000000001"),
    signed("0000101100001011"),
    signed("1110001110101111"),
    signed("0000000000000000"),
    signed("1111110000001001"),
    signed("0010010001011011"),
    signed("0010101010010010"),
    signed("0000001000111001"),
    signed("1111101001100100"),
    signed("0000010101101111"),
    signed("0000010101101111"));

constant lut_gs2q_data_30 : vector_of_signed16(0 to 63) := 
   (signed("1111111011110110"),
    signed("0010010100011100"),
    signed("1111010110100011"),
    signed("1111110101101111"),
    signed("1100110110101001"),
    signed("0000010111010101"),
    signed("0011100100111011"),
    signed("0010100000011111"),
    signed("0000110111100100"),
    signed("0010101010011011"),
    signed("1111101000110101"),
    signed("1101001011100001"),
    signed("1101101011001001"),
    signed("1110100000000011"),
    signed("1111110100111010"),
    signed("1100110101110101"),
    signed("0011010110101101"),
    signed("1110001011010100"),
    signed("0001010111100110"),
    signed("0000010111101001"),
    signed("0011011101010101"),
    signed("0000101011011110"),
    signed("0001110011011111"),
    signed("1100101000111111"),
    signed("0000011111110110"),
    signed("0000111110101000"),
    signed("1101111000100010"),
    signed("1110101011111111"),
    signed("0001110011001010"),
    signed("1111110110110010"),
    signed("1101010011000110"),
    signed("1101011101000001"),
    signed("0001111010010010"),
    signed("1110111011001001"),
    signed("0001000100110111"),
    signed("1101010111100111"),
    signed("0000001011011010"),
    signed("1111111011110001"),
    signed("0000000110110001"),
    signed("1100101001010011"),
    signed("0000001100010010"),
    signed("0001100111011100"),
    signed("1100011010110001"),
    signed("1111101100001101"),
    signed("1111101000000100"),
    signed("0010101101110101"),
    signed("1100110110010101"),
    signed("0010110000001000"),
    signed("1110100100111111"),
    signed("0000011101001100"),
    signed("1110100111000011"),
    signed("0011010111100001"),
    signed("1110101101111101"),
    signed("0011000010101110"),
    signed("0001001100110111"),
    signed("1110001100110110"),
    signed("1111000111100000"),
    signed("0000011100100101"),
    signed("0010011001110110"),
    signed("0010011010101000"),
    signed("1111010000011111"),
    signed("0000010100111111"),
    signed("0001001101011000"),
    signed("0000110111001101"));

constant lut_gs2q_data_31 : vector_of_signed16(0 to 63) := 
   (signed("1111111110111101"),
    signed("0010001111101011"),
    signed("1110100011011111"),
    signed("0000100101010110"),
    signed("1101000100101110"),
    signed("0001001001011000"),
    signed("0011001111101000"),
    signed("0010011011010000"),
    signed("0001101101101111"),
    signed("0010011110100100"),
    signed("1110110010011001"),
    signed("1101001010011000"),
    signed("1101111110001100"),
    signed("1110000011111111"),
    signed("0000011101110000"),
    signed("1100111101001000"),
    signed("0011001010001100"),
    signed("1110010100101001"),
    signed("0001100010100110"),
    signed("0001000111010001"),
    signed("0011001000010101"),
    signed("0001011000100100"),
    signed("0001110100110110"),
    signed("1100110111111011"),
    signed("0000111111000111"),
    signed("0001100000000100"),
    signed("1101111100000011"),
    signed("1110000101010100"),
    signed("0001110110111101"),
    signed("1111010101001111"),
    signed("1101010001101011"),
    signed("1101101100111111"),
    signed("0010010110101001"),
    signed("1110011110101011"),
    signed("0001100001010101"),
    signed("1101011111100011"),
    signed("1111100000001010"),
    signed("0000110101000001"),
    signed("0000111010100001"),
    signed("1100110101110100"),
    signed("1111010110101100"),
    signed("0010001111000110"),
    signed("1100110010011110"),
    signed("1110110100011110"),
    signed("1111000110000110"),
    signed("0010101010001010"),
    signed("1101000110110101"),
    signed("0010101110010001"),
    signed("1110000011111111"),
    signed("0000110111110011"),
    signed("1110000101010100"),
    signed("0011010001110010"),
    signed("1110001011100010"),
    signed("0010111011000101"),
    signed("0001100101100001"),
    signed("1110001001000011"),
    signed("1110010110011100"),
    signed("0001000111010001"),
    signed("0010011101000111"),
    signed("0010001001011010"),
    signed("1110011101111111"),
    signed("0000111111111101"),
    signed("0001111010011111"),
    signed("0001010100100001"));

constant lut_gs2q_data_32 : vector_of_signed16(0 to 63) := 
   (signed("0000000010110111"),
    signed("0010001001011101"),
    signed("1101111100100100"),
    signed("0001010101010111"),
    signed("1101011100111001"),
    signed("0001110100100001"),
    signed("0010101101111001"),
    signed("0010010000010110"),
    signed("0010010100000111"),
    signed("0010001101110000"),
    signed("1110000110000111"),
    signed("1101010100111111"),
    signed("1110001101111010"),
    signed("1101110101010010"),
    signed("0001001001000010"),
    signed("1101010000100101"),
    signed("0010110000110111"),
    signed("1110011000001110"),
    signed("0001110001100010"),
    signed("0001110000110011"),
    signed("0010101000010001"),
    signed("0001111011010101"),
    signed("0001111000100110"),
    signed("1101010010111000"),
    signed("0001011101000101"),
    signed("0001110111110011"),
    signed("1101111110100111"),
    signed("1101101110001100"),
    signed("0001111100010100"),
    signed("1110110001111001"),
    signed("1101011010100111"),
    signed("1101111101001111"),
    signed("0010100000100010"),
    signed("1110001001001011"),
    signed("0001110110110101"),
    signed("1101101101110001"),
    signed("1110110011010000"),
    signed("0001101001101111"),
    signed("0001101001111100"),
    signed("1101001111001001"),
    signed("1110100010100010"),
    signed("0010100011111110"),
    signed("1101010101110110"),
    signed("1110000100100101"),
    signed("1110100100110100"),
    signed("0010011110000110"),
    signed("1101100000101000"),
    signed("0010100010001110"),
    signed("1101110001000110"),
    signed("0001010011010001"),
    signed("1101110010011000"),
    signed("0010111101001011"),
    signed("1101110110000011"),
    signed("0010101000000011"),
    signed("0001110100110101"),
    signed("1110000011101100"),
    signed("1101110011001101"),
    signed("0001101100100110"),
    signed("0010011000111011"),
    signed("0001111010001111"),
    signed("1101111000001010"),
    signed("0001100110111110"),
    signed("0010010110110000"),
    signed("0001101100110100"));

constant lut_gs2q_data_33 : vector_of_signed16(0 to 63) := 
   (signed("0000001001110000"),
    signed("0010000000100101"),
    signed("1101100100100001"),
    signed("0010000000000001"),
    signed("1101111011101001"),
    signed("0010010010111101"),
    signed("0010000000000001"),
    signed("0010000001101101"),
    signed("0010100111011010"),
    signed("0001110110110000"),
    signed("1101100111001011"),
    signed("1101101110101111"),
    signed("1110011001010111"),
    signed("1101110011000111"),
    signed("0001110010000001"),
    signed("1101110001111110"),
    signed("0010001001101011"),
    signed("1110010110101101"),
    signed("0010000000100101"),
    signed("0010001110100111"),
    signed("0001111101010111"),
    signed("0010001101011110"),
    signed("0001111100001110"),
    signed("1101110110010101"),
    signed("0001111011000110"),
    signed("0010000001100011"),
    signed("1101111101010110"),
    signed("1101100111001011"),
    signed("0010000000100101"),
    signed("1110001011111010"),
    signed("1101110001011001"),
    signed("1110001001000110"),
    signed("0010011000110101"),
    signed("1101111000111111"),
    signed("0010000111000001"),
    signed("1110000100010101"),
    signed("1110001001101001"),
    signed("0010010111010011"),
    signed("0010001110100111"),
    signed("1101110001111110"),
    signed("1101110110010101"),
    signed("0010100101001001"),
    signed("1101111111111111"),
    signed("1101100011011001"),
    signed("1110000011001110"),
    signed("0010000111000001"),
    signed("1101111111111111"),
    signed("0010001101101001"),
    signed("1101101100000110"),
    signed("0001101101000101"),
    signed("1101110010100010"),
    signed("0010010111101100"),
    signed("1101101101110011"),
    signed("0010000111100110"),
    signed("0001111100001111"),
    signed("1101111111011011"),
    signed("1101100000001011"),
    signed("0010001011111100"),
    signed("0010001001101011"),
    signed("0001101101101001"),
    signed("1101100001110111"),
    signed("0010000100111100"),
    signed("0010011100000100"),
    signed("0010000001101101"));

constant lut_gs2q_data_34 : vector_of_signed16(0 to 63) := 
   (signed("0000001111001000"),
    signed("0001111000100110"),
    signed("1101100100101000"),
    signed("0010101000101111"),
    signed("1110100101100000"),
    signed("0010100101011001"),
    signed("0001001100000000"),
    signed("0001101000111000"),
    signed("0010100010100111"),
    signed("0001100001000001"),
    signed("1101011111011110"),
    signed("1110010000011100"),
    signed("1110011100011010"),
    signed("1110000100000000"),
    signed("0010011100011010"),
    signed("1110011100111001"),
    signed("0001011001110000"),
    signed("1110001001100000"),
    signed("0010010000100001"),
    signed("0010100101011001"),
    signed("0001001101001110"),
    signed("0010010011010000"),
    signed("0010000101101111"),
    signed("1110100010100010"),
    signed("0010010101011011"),
    signed("0001111110110111"),
    signed("1101111110100111"),
    signed("1101110111011001"),
    signed("0010000101101111"),
    signed("1101100111111100"),
    signed("1110001111001101"),
    signed("1110010001011100"),
    signed("0001111001111001"),
    signed("1101110000101000"),
    signed("0010001111011000"),
    signed("1110011100000101"),
    signed("1101100011100110"),
    signed("0010110011111010"),
    signed("0010101100010000"),
    signed("1110100010100010"),
    signed("1101010010111000"),
    signed("0010001111110001"),
    signed("1110110000010010"),
    signed("1101010000110011"),
    signed("1101101001010111"),
    signed("0001101000001000"),
    signed("1110100101100000"),
    signed("0001101010101101"),
    signed("1101111011111000"),
    signed("0010001010110010"),
    signed("1110000011010000"),
    signed("0001100110000101"),
    signed("1101110110010000"),
    signed("0001100001110100"),
    signed("0001110100110101"),
    signed("1101111010010001"),
    signed("1101100110000100"),
    signed("0010100001000000"),
    signed("0001110001101011"),
    signed("0001100111110010"),
    signed("1101100000011100"),
    signed("0010011110100000"),
    signed("0010001111111010"),
    signed("0010001100011010"));

constant lut_gs2q_data_35 : vector_of_signed16(0 to 63) := 
   (signed("0000010101011001"),
    signed("0001110100110110"),
    signed("1101110110011010"),
    signed("0011000110001110"),
    signed("1111010001010000"),
    signed("0010101110010101"),
    signed("0000011000010011"),
    signed("0001001100111011"),
    signed("0010000100001011"),
    signed("0001000110101101"),
    signed("1101101001010111"),
    signed("1110111110001011"),
    signed("1110010100101001"),
    signed("1110011111111100"),
    signed("0010111110101000"),
    signed("1111001011110000"),
    signed("0000100111001101"),
    signed("1101111000101101"),
    signed("0010100001111011"),
    signed("0010101110010101"),
    signed("0000011101110000"),
    signed("0010000101101000"),
    signed("0010001101100100"),
    signed("1111010110101100"),
    signed("0010101000010001"),
    signed("0001110010010100"),
    signed("1101111100000011"),
    signed("1110010110011100"),
    signed("0010001101100100"),
    signed("1101001010111111"),
    signed("1110111000101111"),
    signed("1110010111111101"),
    signed("0001001101100111"),
    signed("1101110001110011"),
    signed("0010001110001101"),
    signed("1110111010101000"),
    signed("1101000001011000"),
    signed("0011000100110010"),
    signed("0010111011000101"),
    signed("1111010110101100"),
    signed("1100110111111011"),
    signed("0001100100001000"),
    signed("1111100101100110"),
    signed("1101001010011000"),
    signed("1101010010010011"),
    signed("0001000101011000"),
    signed("1111010001010000"),
    signed("0001000010000100"),
    signed("1110011000010101"),
    signed("0010100100000000"),
    signed("1110100000001001"),
    signed("0000101110110100"),
    signed("1110010001000010"),
    signed("0000110010111011"),
    signed("0001100101100001"),
    signed("1101110010011100"),
    signed("1101111101101110"),
    signed("0010101000110101"),
    signed("0001010100010010"),
    signed("0001101011010111"),
    signed("1101110110011010"),
    signed("0010101100001011"),
    signed("0001101101101111"),
    signed("0010010011101010"));

constant lut_gs2q_data_36 : vector_of_signed16(0 to 63) := 
   (signed("0000011101001101"),
    signed("0001110011011111"),
    signed("1110011001101101"),
    signed("0011011000101110"),
    signed("1111111110000100"),
    signed("0010101100111010"),
    signed("1111100110101100"),
    signed("0000101100100001"),
    signed("0001010010110100"),
    signed("0000101010100010"),
    signed("1110000101101110"),
    signed("1111110001101001"),
    signed("1110000110011001"),
    signed("1111000110010011"),
    signed("0011010111111001"),
    signed("1111111100111011"),
    signed("1111110100000010"),
    signed("1101100101000100"),
    signed("0010110000010101"),
    signed("0010101100111010"),
    signed("1111101111111111"),
    signed("0001101000010100"),
    signed("0010010100110001"),
    signed("0000001100010010"),
    signed("0010110100110010"),
    signed("0001011010100001"),
    signed("1101111000100010"),
    signed("1111000010100101"),
    signed("0010010100110001"),
    signed("1100110101011010"),
    signed("1111101000010111"),
    signed("1110011010001100"),
    signed("0000010111001011"),
    signed("1101111000011011"),
    signed("0010000111100101"),
    signed("1111011100011110"),
    signed("1100101000000111"),
    signed("0011001000001010"),
    signed("0010111101110010"),
    signed("0000001100010010"),
    signed("1100101000111111"),
    signed("0000101010010001"),
    signed("0000011001101000"),
    signed("1101010000011100"),
    signed("1101000001111011"),
    signed("0000011110100111"),
    signed("1111111110000100"),
    signed("0000010100101011"),
    signed("1111000000100011"),
    signed("0010111000101001"),
    signed("1111001000000000"),
    signed("1111110100110111"),
    signed("1110111000111101"),
    signed("0000000001000001"),
    signed("0001001100110111"),
    signed("1101101011001111"),
    signed("1110100110001110"),
    signed("0010100110110101"),
    signed("0000110000111000"),
    signed("0001110100101100"),
    signed("1110011110101001"),
    signed("0010110000011100"),
    signed("0000111100100000"),
    signed("0010010101110011"));

constant lut_gs2q_data_37 : vector_of_signed16(0 to 63) := 
   (signed("0000100111010110"),
    signed("0001110100011001"),
    signed("1111001010000111"),
    signed("0011011111000001"),
    signed("0000101000101110"),
    signed("0010100011101101"),
    signed("1110111010111110"),
    signed("0000001000111001"),
    signed("0000010101101111"),
    signed("0000001100110110"),
    signed("1110110001010000"),
    signed("0000100101100110"),
    signed("1101110101001010"),
    signed("1111110011010001"),
    signed("0011100101100111"),
    signed("0000101100001011"),
    signed("1111000100101011"),
    signed("1101010010100110"),
    signed("0010111001011100"),
    signed("0010100011101101"),
    signed("1111000110111111"),
    signed("0000111110011101"),
    signed("0010011001111111"),
    signed("0000111110011101"),
    signed("0010111010001001"),
    signed("0000111001000001"),
    signed("1101110101001010"),
    signed("1111110110010010"),
    signed("0010011001111111"),
    signed("1100101001100011"),
    signed("0000011001100100"),
    signed("1110011000011100"),
    signed("1111011101011011"),
    signed("1110000010000000"),
    signed("0001111110000000"),
    signed("0000000000000000"),
    signed("1100011010011001"),
    signed("0011000000000001"),
    signed("0010110110010100"),
    signed("0000111110011101"),
    signed("1100100110011011"),
    signed("1111101010010001"),
    signed("0001001000001010"),
    signed("1101011111011011"),
    signed("1100111001110110"),
    signed("1111110110010010"),
    signed("0000101000101110"),
    signed("1111100110011100"),
    signed("1111110000001001"),
    signed("0011000110001010"),
    signed("1111110110010010"),
    signed("1110111110000110"),
    signed("1111101001100100"),
    signed("1111010000101101"),
    signed("0000101100001011"),
    signed("1101100110000001"),
    signed("1111011010011010"),
    signed("0010011101011101"),
    signed("0000001001101110"),
    signed("0010000001001000"),
    signed("1111010011110101"),
    signed("0010101100100110"),
    signed("0000000011001000"),
    signed("0010010011101111"));

constant lut_gs2q_data_38 : vector_of_signed16(0 to 63) := 
   (signed("0000110100101001"),
    signed("0001110111001011"),
    signed("0000000001110101"),
    signed("0011011000101110"),
    signed("0001001110000000"),
    signed("0010010110000000"),
    signed("1110011000100000"),
    signed("1111100011101100"),
    signed("1111010101101111"),
    signed("1111101101110100"),
    signed("1111100111001100"),
    signed("0001010100010110"),
    signed("1101100101010101"),
    signed("0000100010010101"),
    signed("0011100101110000"),
    signed("0001010101010001"),
    signed("1110011101011100"),
    signed("1101000101110000"),
    signed("0010111011001000"),
    signed("0010010110000000"),
    signed("1110100101011111"),
    signed("0000001100010010"),
    signed("0010011011111000"),
    signed("0001101000010100"),
    signed("0010110111110001"),
    signed("0000010000000001"),
    signed("1101110011001011"),
    signed("0000101011001010"),
    signed("0010011011111000"),
    signed("1100101001010011"),
    signed("0001000111010111"),
    signed("1110010011100001"),
    signed("1110100111111100"),
    signed("1110001011101001"),
    signed("0001110100010111"),
    signed("0000100011100010"),
    signed("1100011010010000"),
    signed("0010101111100000"),
    signed("0010100111100110"),
    signed("0001101000010100"),
    signed("1100101111101001"),
    signed("1110101101001100"),
    signed("0001101101010000"),
    signed("1101110010101110"),
    signed("1100111011010001"),
    signed("1111001111001000"),
    signed("0001001110000000"),
    signed("1110111011100111"),
    signed("0000100010000001"),
    signed("0011001010001011"),
    signed("0000100101101110"),
    signed("1110010000011010"),
    signed("0000011101011010"),
    signed("1110100110101111"),
    signed("0000000101010101"),
    signed("1101100100001000"),
    signed("0000010011110011"),
    signed("0010001111111100"),
    signed("1111100001011001"),
    signed("0010001101010101"),
    signed("0000001111001011"),
    signed("0010100010101010"),
    signed("1111001001100101"),
    signed("0010001110101100"));

constant lut_gs2q_data_39 : vector_of_signed16(0 to 63) := 
   (signed("0001000101100110"),
    signed("0001111011000111"),
    signed("0000111010100001"),
    signed("0011000110001110"),
    signed("0001101011000001"),
    signed("0010000111010011"),
    signed("1110000001111110"),
    signed("1110111110101111"),
    signed("1110011011111000"),
    signed("1111001101101101"),
    signed("0000100010000000"),
    signed("0001111000100101"),
    signed("1101011011010010"),
    signed("0001001110111000"),
    signed("0011010111001111"),
    signed("0001110100011011"),
    signed("1110000001111110"),
    signed("1101000010110001"),
    signed("0010110011110001"),
    signed("0010000111010011"),
    signed("1110001101101100"),
    signed("1111010110101100"),
    signed("0010011001001010"),
    signed("0010000101101000"),
    signed("0010101101011110"),
    signed("1111100010010000"),
    signed("1101110011111001"),
    signed("0001011010101010"),
    signed("0010011001001010"),
    signed("1100110101110100"),
    signed("0001101100111000"),
    signed("1110001100011111"),
    signed("1101111101111011"),
    signed("1110010010100011"),
    signed("0001101101011101"),
    signed("0001000101011000"),
    signed("1100101000110001"),
    signed("0010011010010100"),
    signed("0010010101000111"),
    signed("0010000101101000"),
    signed("1101000011011001"),
    signed("1101111011110101"),
    signed("0010000101101000"),
    signed("1110000101100000"),
    signed("1101000110110101"),
    signed("1110101011101110"),
    signed("0001101011000001"),
    signed("1110011000010101"),
    signed("0001010000111110"),
    signed("0011000010111000"),
    signed("0001010000111101"),
    signed("1101110000111110"),
    signed("0001001110111000"),
    signed("1110000111011011"),
    signed("1111011010101010"),
    signed("1101100110110110"),
    signed("0001001011100010"),
    signed("0010000001110100"),
    signed("1110111010101000"),
    signed("0010010101110100"),
    signed("0001001001011011"),
    signed("0010010101000111"),
    signed("1110010111110001"),
    signed("0010001000000100"));

constant lut_gs2q_data_40 : vector_of_signed16(0 to 63) := 
   (signed("0001011010010001"),
    signed("0001111111011011"),
    signed("0001101110001001"),
    signed("0010101000101111"),
    signed("0001111101011100"),
    signed("0001111010101101"),
    signed("1101111001000101"),
    signed("1110011100000001"),
    signed("1101110000001111"),
    signed("1110101100111100"),
    signed("0001011100000011"),
    signed("0010001110000101"),
    signed("1101011010110000"),
    signed("0001110100101110"),
    signed("0010111010001101"),
    signed("0010000110110010"),
    signed("1101110100111001"),
    signed("1101001100110111"),
    signed("0010100010011011"),
    signed("0001111010101101"),
    signed("1110000001001001"),
    signed("1110100010100010"),
    signed("0010010000110100"),
    signed("0010010011010000"),
    signed("0010011011100000"),
    signed("1110110010110010"),
    signed("1101111000100011"),
    signed("0001111111000011"),
    signed("0010010000110100"),
    signed("1101001111001001"),
    signed("0010000110000001"),
    signed("1110000100100000"),
    signed("1101100101010100"),
    signed("1110010100011111"),
    signed("0001101011100001"),
    signed("0001100011111011"),
    signed("1101000101110011"),
    signed("0010000100001100"),
    signed("0010000010010011"),
    signed("0010010011010000"),
    signed("1101011111110011"),
    signed("1101011101011001"),
    signed("0010001111000011"),
    signed("1110010011100001"),
    signed("1101011100011011"),
    signed("1110001110010101"),
    signed("0001111101011100"),
    signed("1110000000000100"),
    signed("0001111000011101"),
    signed("0010101111011011"),
    signed("0001110011001100"),
    signed("1101100011011010"),
    signed("0001111000111011"),
    signed("1101110110000111"),
    signed("1110101110110110"),
    signed("1101101111001100"),
    signed("0001111011011011"),
    signed("0001110110010011"),
    signed("1110010111111000"),
    signed("0010010111100000"),
    signed("0001111011111001"),
    signed("0010000110011111"),
    signed("1101110100011111"),
    signed("0010000001010101"));

constant lut_gs2q_data_41 : vector_of_signed16(0 to 63) := 
   (signed("0001110100001011"),
    signed("0010000101100000"),
    signed("0010010101100111"),
    signed("0010000000000001"),
    signed("0010000001100011"),
    signed("0001110100101001"),
    signed("1101111100001100"),
    signed("1101111011010000"),
    signed("1101011010110111"),
    signed("1110001110100100"),
    signed("0010010010011000"),
    signed("0010010000001000"),
    signed("1101100011111110"),
    signed("0010001110100111"),
    signed("0010001110000010"),
    signed("0010001100111001"),
    signed("1101110101001100"),
    signed("1101100011011001"),
    signed("0010000100111100"),
    signed("0001110100101001"),
    signed("1101111110011101"),
    signed("1101110001111110"),
    signed("0010000000000001"),
    signed("0010010001110100"),
    signed("0010000100110000"),
    signed("1110000010101001"),
    signed("1101111111111111"),
    signed("0010010001110100"),
    signed("0010000000000001"),
    signed("1101110110010101"),
    signed("0010001101110111"),
    signed("1101111110110110"),
    signed("1101011111100110"),
    signed("1110010010010111"),
    signed("0001110001111111"),
    signed("0010000000000001"),
    signed("1101101101101000"),
    signed("0001101110001110"),
    signed("0001101111111010"),
    signed("0010010001110100"),
    signed("1110000100111010"),
    signed("1101010100010000"),
    signed("0010001010110100"),
    signed("1110010111101011"),
    signed("1101111000111111"),
    signed("1101110110010101"),
    signed("0010000001100011"),
    signed("1101110011000111"),
    signed("0010010111010011"),
    signed("0010001110000010"),
    signed("0010001010110100"),
    signed("1101100111001011"),
    signed("0010010101100111"),
    signed("1101110110111000"),
    signed("1110000110111111"),
    signed("1101111111111111"),
    signed("0010011100100111"),
    signed("0001101101101001"),
    signed("1101111101010101"),
    signed("0010010010011000"),
    signed("0010011111010001"),
    signed("0001110110111010"),
    signed("1101100110100110"),
    signed("0001111001100100"));

constant lut_gs2q_data_42 : vector_of_signed16(0 to 63) := 
   (signed("0010001101001100"),
    signed("0010001010000000"),
    signed("0010110100011000"),
    signed("0001010101010111"),
    signed("0001111101011100"),
    signed("0001110011101001"),
    signed("1110001101010010"),
    signed("1101100000110001"),
    signed("1101011100000010"),
    signed("1101110001010010"),
    signed("0010111010001101"),
    signed("0010000100111000"),
    signed("1101111110010010"),
    signed("0010100001011110"),
    signed("0001011000010101"),
    signed("0001111111111100"),
    signed("1110000101001001"),
    signed("1110001000100001"),
    signed("0001100011000011"),
    signed("0001110011101001"),
    signed("1110001000001101"),
    signed("1101001111001001"),
    signed("0001101101010010"),
    signed("0001111111000011"),
    signed("0001100111101110"),
    signed("1101010111101111"),
    signed("1110001101100100"),
    signed("0010010011010000"),
    signed("0001101101010010"),
    signed("1110100110010000"),
    signed("0010001001111101"),
    signed("1101110101110011"),
    signed("1101110000010011"),
    signed("1110001001100000"),
    signed("0001111010001111"),
    signed("0010010101111101"),
    signed("1110100011111101"),
    signed("0001100001011111"),
    signed("0001100010101101"),
    signed("0001111111000011"),
    signed("1110101101101101"),
    signed("1101101000001011"),
    signed("0001110110111011"),
    signed("1110010111011101"),
    signed("1110011101010111"),
    signed("1101100111000101"),
    signed("0001111101011100"),
    signed("1101111001001110"),
    signed("0010100101001100"),
    signed("0001100011000111"),
    signed("0010010010110010"),
    signed("1110000010001011"),
    signed("0010101001100110"),
    signed("1110000011010000"),
    signed("1101011111011001"),
    signed("1110010010101110"),
    signed("0010101111001101"),
    signed("0001101011101110"),
    signed("1101100101101001"),
    signed("0001111110110000"),
    signed("0010110111010110"),
    signed("0001101010110110"),
    signed("1101101101011100"),
    signed("0001110100011001"));

constant lut_gs2q_data_43 : vector_of_signed16(0 to 63) := 
   (signed("0010100101000100"),
    signed("0010001001111110"),
    signed("0011000010101011"),
    signed("0000100101010110"),
    signed("0001101011000001"),
    signed("0001110101000011"),
    signed("1110101100111100"),
    signed("1101010000011011"),
    signed("1101110000111010"),
    signed("1101010100011001"),
    signed("0011010111001111"),
    signed("0001100111011110"),
    signed("1110100010000001"),
    signed("0010100110101110"),
    signed("0000011111111010"),
    signed("0001100111101011"),
    signed("1110100101010110"),
    signed("1110111100000101"),
    signed("0000111000010111"),
    signed("0001110101000011"),
    signed("1110011111111100"),
    signed("1100110101110100"),
    signed("0001010010011011"),
    signed("0001011010101010"),
    signed("0001000011010111"),
    signed("1100110111101011"),
    signed("1110100100001011"),
    signed("0010000101101000"),
    signed("0001010010011011"),
    signed("1111011000110011"),
    signed("0001110100011110"),
    signed("1101110000100010"),
    signed("1110010111110001"),
    signed("1101111000101101"),
    signed("0010001001011010"),
    signed("0010100010100100"),
    signed("1111011110000000"),
    signed("0001011000111001"),
    signed("0001011110010110"),
    signed("0001011010101010"),
    signed("1111010101001111"),
    signed("1110010000001011"),
    signed("0001010011000100"),
    signed("1110001101000110"),
    signed("1111001001101001"),
    signed("1101100010111001"),
    signed("0001101011000001"),
    signed("1110001011100101"),
    signed("0010101000110101"),
    signed("0000110100010000"),
    signed("0010000111101111"),
    signed("1110101010110010"),
    signed("0010101110010101"),
    signed("1110100000001001"),
    signed("1101000001011000"),
    signed("1110101101100101"),
    signed("0010110101101000"),
    signed("0001110010111101"),
    signed("1101010111111100"),
    signed("0001100011011011"),
    signed("0010111101001111"),
    signed("0001100101111100"),
    signed("1110000101100001"),
    signed("0001110100110110"));

constant lut_gs2q_data_44 : vector_of_signed16(0 to 63) := 
   (signed("0010111001000110"),
    signed("0010000111101111"),
    signed("0011000011100010"),
    signed("1111110101101111"),
    signed("0001001110000000"),
    signed("0001111010001000"),
    signed("1111010101101011"),
    signed("1101001000100100"),
    signed("1110011000100100"),
    signed("1100111100101011"),
    signed("0011100101110000"),
    signed("0000111101110000"),
    signed("1111001110100111"),
    signed("0010100010001110"),
    signed("1111100111100001"),
    signed("0001000100011001"),
    signed("1111001111111011"),
    signed("1111110110111001"),
    signed("0000001010010011"),
    signed("0001111010001000"),
    signed("1111000001011000"),
    signed("1100101001010011"),
    signed("0000110010100101"),
    signed("0000101011001010"),
    signed("0000011100000000"),
    signed("1100100010101011"),
    signed("1111000001001110"),
    signed("0001101000010100"),
    signed("0000110010100101"),
    signed("0000001011111110"),
    signed("0001010010000011"),
    signed("1101101101010001"),
    signed("1111001110100000"),
    signed("1101100101000100"),
    signed("0010011010101000"),
    signed("0010101000000101"),
    signed("0000011000110100"),
    signed("0001010111000110"),
    signed("0001100000011000"),
    signed("0000101011001010"),
    signed("1111111011101110"),
    signed("1111001000110000"),
    signed("0000100101011001"),
    signed("1101111101011010"),
    signed("1111111000010100"),
    signed("1101100110001010"),
    signed("0001001110000000"),
    signed("1110101010101111"),
    signed("0010100001111001"),
    signed("0000000011000101"),
    signed("0001101100111100"),
    signed("1111011110001001"),
    signed("0010100111111110"),
    signed("1111001000000000"),
    signed("1100101101000010"),
    signed("1111001101011011"),
    signed("0010101111100100"),
    signed("0001111111011000"),
    signed("1101010001110111"),
    signed("0000111111100111"),
    signed("0010110101010100"),
    signed("0001100110001001"),
    signed("1110101101101100"),
    signed("0001111000011010"));

constant lut_gs2q_data_45 : vector_of_signed16(0 to 63) := 
   (signed("0011000110011001"),
    signed("0010000011111000"),
    signed("0010111001011100"),
    signed("1111001010000111"),
    signed("0000101000101110"),
    signed("0010000001001000"),
    signed("0000000011001000"),
    signed("1101001000111111"),
    signed("1111001101100101"),
    signed("1100101101000000"),
    signed("0011100101100111"),
    signed("0000001100110110"),
    signed("0000000000000000"),
    signed("0010010110110111"),
    signed("1110110100011000"),
    signed("0000011001100100"),
    signed("0000000000000000"),
    signed("0000110010011011"),
    signed("1111011100101110"),
    signed("0010000001001000"),
    signed("1111101001100100"),
    signed("1100101001100011"),
    signed("0000001111001001"),
    signed("1111110110010010"),
    signed("1111110011111111"),
    signed("1100011010011001"),
    signed("1111100011101011"),
    signed("0000111110011101"),
    signed("0000001111001001"),
    signed("0000111011010101"),
    signed("0000100110011010"),
    signed("1101101100001010"),
    signed("0000001100110110"),
    signed("1101010010100110"),
    signed("0010101010010010"),
    signed("0010100111001010"),
    signed("0001001110110000"),
    signed("0001011011100010"),
    signed("0001100111100100"),
    signed("1111110110010010"),
    signed("0000011111011101"),
    signed("0000001001101110"),
    signed("1111110011001010"),
    signed("1101101100010001"),
    signed("0000100101100110"),
    signed("1101101110100101"),
    signed("0000101000101110"),
    signed("1111010011110101"),
    signed("0010010011101111"),
    signed("1111010011110101"),
    signed("0001000101000010"),
    signed("0000010101101111"),
    signed("0010011001111111"),
    signed("1111110110010010"),
    signed("1100100100000111"),
    signed("1111110000110111"),
    signed("0010100000100101"),
    signed("0010001101111110"),
    signed("1101010010100110"),
    signed("0000010101101111"),
    signed("0010100011101101"),
    signed("0001101010101100"),
    signed("1111100000100011"),
    signed("0001111110000111"));

constant lut_gs2q_data_46 : vector_of_signed16(0 to 63) := 
   (signed("0011001010001111"),
    signed("0001111111010100"),
    signed("0010100111111011"),
    signed("1110100101110011"),
    signed("1111111110000100"),
    signed("0010000111111001"),
    signed("0000110000011010"),
    signed("1101010000111110"),
    signed("0000001001000111"),
    signed("1100101000001010"),
    signed("0011010111111001"),
    signed("1111011010100111"),
    signed("0000110001011001"),
    signed("0010001000010110"),
    signed("1110001011011111"),
    signed("1111101011010101"),
    signed("0000110000000101"),
    signed("0001100111011100"),
    signed("1110110011101101"),
    signed("0010000111111001"),
    signed("0000010100111111"),
    signed("1100110101011010"),
    signed("1111101001110001"),
    signed("1111000010100101"),
    signed("1111001101101111"),
    signed("1100011111101100"),
    signed("0000001010000010"),
    signed("0000001100010010"),
    signed("1111101001110001"),
    signed("0001100010100100"),
    signed("1111110110000001"),
    signed("1101101101010001"),
    signed("0001001001110110"),
    signed("1101000101110000"),
    signed("0010110100011111"),
    signed("0010100000111110"),
    signed("0001111010010010"),
    signed("0001100100111100"),
    signed("0001110001111010"),
    signed("1111000010100101"),
    signed("0000111111000111"),
    signed("0001001001100010"),
    signed("1111000010010000"),
    signed("1101011110000111"),
    signed("0001001101101011"),
    signed("1101111001010111"),
    signed("1111111110000100"),
    signed("0000000011000101"),
    signed("0010000010100110"),
    signed("1110101010101111"),
    signed("0000010011111000"),
    signed("0001001010011010"),
    signed("0010001000101010"),
    signed("0000100101101110"),
    signed("1100100111100111"),
    signed("0000010110001111"),
    signed("0010001101010010"),
    signed("0010011010111111"),
    signed("1101011000111110"),
    signed("1111101000111100"),
    signed("0010001101100110"),
    signed("0001110010001111"),
    signed("0000010111100000"),
    signed("0010000100100001"));

constant lut_gs2q_data_47 : vector_of_signed16(0 to 63) := 
   (signed("0011000010101000"),
    signed("0001111011000100"),
    signed("0010010011000001"),
    signed("1110001011100101"),
    signed("1111010001010000"),
    signed("0010001100000111"),
    signed("0001011000100100"),
    signed("1101011111010101"),
    signed("0001000011111011"),
    signed("1100110000010100"),
    signed("0010111110101000"),
    signed("1110101100111100"),
    signed("0001011101111111"),
    signed("0001111010100000"),
    signed("1101110000111110"),
    signed("1110111101111100"),
    signed("0001011010101010"),
    signed("0010001111000110"),
    signed("1110010011001000"),
    signed("0010001100000111"),
    signed("0000111111111101"),
    signed("1101001010111111"),
    signed("1111000100001111"),
    signed("1110010110011100"),
    signed("1110101011011111"),
    signed("1100110010011110"),
    signed("0000110010010111"),
    signed("1111010110101100"),
    signed("1111000100001111"),
    signed("0001111110000010"),
    signed("1111000101100010"),
    signed("1101110000100010"),
    signed("0001111100101001"),
    signed("1101000010110001"),
    signed("0010110101101000"),
    signed("0010010110111110"),
    signed("0010010110101001"),
    signed("0001110001100000"),
    signed("0001111101001110"),
    signed("1110010110011100"),
    signed("0001011001101110"),
    signed("0001111110101111"),
    signed("1110011000100010"),
    signed("1101010111001011"),
    signed("0001101101000111"),
    signed("1110000011101001"),
    signed("1111010001010000"),
    signed("0000110100010000"),
    signed("0001110010111010"),
    signed("1110001011100101"),
    signed("1111011110000000"),
    signed("0001110101010001"),
    signed("0001111000011001"),
    signed("0001010000111101"),
    signed("1100110111101011"),
    signed("0000111011110001"),
    signed("0001111010100000"),
    signed("0010100010100111"),
    signed("1101100011100010"),
    signed("1110111100101001"),
    signed("0001111000011001"),
    signed("0001111011000111"),
    signed("0001001011100001"),
    signed("0010001010000001"));

constant lut_gs2q_data_48 : vector_of_signed16(0 to 63) := 
   (signed("0010101110100011"),
    signed("0001111000000100"),
    signed("0001111110100100"),
    signed("1101111101011011"),
    signed("1110100101100000"),
    signed("0010001011101001"),
    signed("0001110111001000"),
    signed("1101110010101110"),
    signed("0001110111011111"),
    signed("1101000110100011"),
    signed("0010011100011010"),
    signed("1110001001000101"),
    signed("0010000001101110"),
    signed("0001110000101011"),
    signed("1101100111100110"),
    signed("1110010101010011"),
    signed("0001111010110111"),
    signed("0010100011111110"),
    signed("1101111110001011"),
    signed("0010001011101001"),
    signed("0001100110111110"),
    signed("1101100111111100"),
    signed("1110100000011011"),
    signed("1101110111011001"),
    signed("1110001111000000"),
    signed("1101010001101001"),
    signed("0001011010011100"),
    signed("1110100010100010"),
    signed("1110100000011011"),
    signed("0010001011000111"),
    signed("1110011001001111"),
    signed("1101110101110011"),
    signed("0010011101101010"),
    signed("1101001100110111"),
    signed("0010101011000001"),
    signed("0010001010111001"),
    signed("0010100000100010"),
    signed("0001111111010010"),
    signed("0010000111010110"),
    signed("1101110111011001"),
    signed("0001101110101101"),
    signed("0010100001011001"),
    signed("1101111011001000"),
    signed("1101011010110100"),
    signed("0010000001001010"),
    signed("1110001010111100"),
    signed("1110100101100000"),
    signed("0001100011000111"),
    signed("0001101000100011"),
    signed("1101111001001110"),
    signed("1110101000001001"),
    signed("0010010000101011"),
    signed("0001101100111101"),
    signed("0001110011001100"),
    signed("1101010011100011"),
    signed("0001011111100101"),
    signed("0001101100011111"),
    signed("0010100001100010"),
    signed("1101110000101110"),
    signed("1110010100000110"),
    signed("0001101000110000"),
    signed("0010000011101000"),
    signed("0001110110001010"),
    signed("0010001101001011"));

constant lut_gs2q_data_49 : vector_of_signed16(0 to 63) := 
   (signed("0010001100001001"),
    signed("0001110100110101"),
    signed("0001101111111010"),
    signed("1101111110011101"),
    signed("1101111111111111"),
    signed("0010000010101011"),
    signed("0010000110011110"),
    signed("1110001011111010"),
    signed("0010011100100111"),
    signed("1101101000010100"),
    signed("0001110110010111"),
    signed("1101110101001100"),
    signed("0010010111101100"),
    signed("0001101111010101"),
    signed("1101110010100010"),
    signed("1101110010010111"),
    signed("0010001111001010"),
    signed("0010100000110011"),
    signed("1101111001001001"),
    signed("0010000010101011"),
    signed("0010001001010010"),
    signed("1110000111100100"),
    signed("1110000010010000"),
    signed("1101101011100010"),
    signed("1101111011101001"),
    signed("1101111101010101"),
    signed("0001111101110000"),
    signed("1101110001111110"),
    signed("1101111101111010"),
    signed("0010001010110100"),
    signed("1101110110101110"),
    signed("1101111110110110"),
    signed("0010100101101110"),
    signed("1101100111101111"),
    signed("0010010101100111"),
    signed("0001111100001110"),
    signed("0010011000110101"),
    signed("0010001110100101"),
    signed("0010010000110110"),
    signed("1101100111001011"),
    signed("0010000000000001"),
    signed("0010101110011010"),
    signed("1101101011100010"),
    signed("1101101000101101"),
    signed("0010000101111001"),
    signed("1110001111101101"),
    signed("1101111011101001"),
    signed("0010001001101011"),
    signed("0001101000010101"),
    signed("1101110011000111"),
    signed("1101110100101000"),
    signed("0010010110110000"),
    signed("0001100110101001"),
    signed("0010001010110100"),
    signed("1101111011101001"),
    signed("0001111101110000"),
    signed("0001101000010101"),
    signed("0010010011010110"),
    signed("1101111100110001"),
    signed("1101101111111001"),
    signed("0001100011111111"),
    signed("0010001100100000"),
    signed("0010010100011110"),
    signed("0010001111001010"));

constant lut_gs2q_data_50 : vector_of_signed16(0 to 63) := 
   (signed("0001100001110110"),
    signed("0001110100010101"),
    signed("0001100110011100"),
    signed("1110001011111011"),
    signed("1101100000101000"),
    signed("0001110110110101"),
    signed("0010001011000111"),
    signed("1110100111000111"),
    signed("0010110011001001"),
    signed("1110010110001101"),
    signed("0001001100110000"),
    signed("1101110000111101"),
    signed("0010100001100010"),
    signed("0001110000101011"),
    signed("1110001110000010"),
    signed("1101011101110010"),
    signed("0010001110110110"),
    signed("0010001100000011"),
    signed("1101111110001011"),
    signed("0001110110110101"),
    signed("0010100010001110"),
    signed("1110101110001011"),
    signed("1101101000101100"),
    signed("1101110001111011"),
    signed("1101101111001100"),
    signed("1110101011111000"),
    signed("0010100000101011"),
    signed("1101001111001001"),
    signed("1101100100111110"),
    signed("0001111010110111"),
    signed("1101011101100101"),
    signed("1110000100100000"),
    signed("0010011001101110"),
    signed("1110001100001111"),
    signed("0001110011010011"),
    signed("0001101111001111"),
    signed("0001111001111001"),
    signed("0010010111001101"),
    signed("0010010010001000"),
    signed("1101101110001100"),
    signed("0010001011001011"),
    signed("0010011101011101"),
    signed("1101101110001100"),
    signed("1110000111100011"),
    signed("0001111101011100"),
    signed("1110001110101010"),
    signed("1101011100111001"),
    signed("0010101011101101"),
    signed("0001101100011111"),
    signed("1110000000000100"),
    signed("1101001101111011"),
    signed("0010001001000000"),
    signed("0001101100111101"),
    signed("0010010010110010"),
    signed("1110101010101001"),
    signed("0010010111010100"),
    signed("0001101000100011"),
    signed("0001111110000000"),
    signed("1110001000110110"),
    signed("1101011000101001"),
    signed("0001101000100011"),
    signed("0010010010001000"),
    signed("0010100000100010"),
    signed("0010001100111110"));

constant lut_gs2q_data_51 : vector_of_signed16(0 to 63) := 
   (signed("0000110000110111"),
    signed("0001111000111101"),
    signed("0001100000011100"),
    signed("1110100010000010"),
    signed("1101000110110101"),
    signed("0001100001010101"),
    signed("0001111110000010"),
    signed("1111000000111001"),
    signed("0010111101001111"),
    signed("1111001111000110"),
    signed("0000011111110110"),
    signed("1101111010011000"),
    signed("0010100010100111"),
    signed("0001111010100000"),
    signed("1110110100011111"),
    signed("1101010001101111"),
    signed("0010000000001000"),
    signed("0001100010000001"),
    signed("1110010011001000"),
    signed("0001100001010101"),
    signed("0010101110010001"),
    signed("1111010011001001"),
    signed("1101010010100010"),
    signed("1110000111011011"),
    signed("1101100110110110"),
    signed("1111100000000110"),
    signed("0010111010100001"),
    signed("1100110101110100"),
    signed("1101010000011011"),
    signed("0001011010101010"),
    signed("1101001100001111"),
    signed("1110001100011111"),
    signed("0001110101000010"),
    signed("1110111110001011"),
    signed("0001000011111011"),
    signed("0001100111110011"),
    signed("0001001101100111"),
    signed("0010011110100101"),
    signed("0010010001100100"),
    signed("1110000101010100"),
    signed("0010001110001101"),
    signed("0001110111001001"),
    signed("1110000101010100"),
    signed("1110101111000010"),
    signed("0001101011000001"),
    signed("1110000101101111"),
    signed("1101000100101110"),
    signed("0011000000110010"),
    signed("0001111010100000"),
    signed("1110011000010101"),
    signed("1100110000011000"),
    signed("0001101011100101"),
    signed("0001111000011001"),
    signed("0010000111101111"),
    signed("1111011010101010"),
    signed("0010101101011110"),
    signed("0001110010111010"),
    signed("0001011011111000"),
    signed("1110010110000110"),
    signed("1101001000110101"),
    signed("0001110010111010"),
    signed("0010010001100100"),
    signed("0010010110101001"),
    signed("0010000100100001"));

constant lut_gs2q_data_52 : vector_of_signed16(0 to 63) := 
   (signed("1111111101011010"),
    signed("0001111111101001"),
    signed("0001100000000100"),
    signed("1111000001000011"),
    signed("1100110110010101"),
    signed("0001000100110111"),
    signed("0001100010100100"),
    signed("1111011011001110"),
    signed("0010111010010000"),
    signed("0000001011011110"),
    signed("1111110100100110"),
    signed("1110010010110000"),
    signed("0010011010111111"),
    signed("0010001000010110"),
    signed("1111100011100101"),
    signed("1101001111111000"),
    signed("0001100010010000"),
    signed("0000101010100110"),
    signed("1110110011101101"),
    signed("0001000100110111"),
    signed("0010110000001000"),
    signed("1111110111000111"),
    signed("1101000011010100"),
    signed("1110101011101010"),
    signed("1101100100001000"),
    signed("0000010011100100"),
    signed("0011001011101111"),
    signed("1100101001010011"),
    signed("1101000011101000"),
    signed("0000110000000101"),
    signed("1101000100111000"),
    signed("1110010011100001"),
    signed("0000111111001010"),
    signed("1111110110100101"),
    signed("0000001110000010"),
    signed("0001100100011100"),
    signed("0000010111001011"),
    signed("0010100001110010"),
    signed("0010001101011111"),
    signed("1110101011111111"),
    signed("0010001100100000"),
    signed("0000111110110110"),
    signed("1110101011111111"),
    signed("1111011101111111"),
    signed("0001001110000000"),
    signed("1101111001000011"),
    signed("1100110110101001"),
    signed("0011001010100000"),
    signed("0010001101010010"),
    signed("1110111011100111"),
    signed("1100100000000001"),
    signed("0001000000000010"),
    signed("0010001000101010"),
    signed("0001101100111100"),
    signed("0000001010010001"),
    signed("0010111100101100"),
    signed("0010000010100110"),
    signed("0000110001101101"),
    signed("1110100000110100"),
    signed("1101000010110011"),
    signed("0010000010100110"),
    signed("0010001101011111"),
    signed("0001111010010010"),
    signed("0001111001100000"));

constant lut_gs2q_data_53 : vector_of_signed16(0 to 63) := 
   (signed("1111001100010000"),
    signed("0010000111000000"),
    signed("0001100100011100"),
    signed("1111100110011100"),
    signed("1100110000001000"),
    signed("0000100010100101"),
    signed("0000111011010101"),
    signed("1111110110010010"),
    signed("0010101101011010"),
    signed("0001000101000010"),
    signed("1111001101100101"),
    signed("1110110111110110"),
    signed("0010001101111110"),
    signed("0010010110110111"),
    signed("0000010101101111"),
    signed("1101010110100010"),
    signed("0000111000001101"),
    signed("1111101101011001"),
    signed("1111011100101110"),
    signed("0000100010100101"),
    signed("0010101001011110"),
    signed("0000011000110111"),
    signed("1100111100001010"),
    signed("1111011010011010"),
    signed("1101100110000001"),
    signed("0001000001111010"),
    signed("0011010011000000"),
    signed("1100101001100011"),
    signed("1100111111010010"),
    signed("0000000000000000"),
    signed("1101000110100100"),
    signed("1110011000011100"),
    signed("0000000000000000"),
    signed("0000101111010011"),
    signed("1111010111010010"),
    signed("0001100101010000"),
    signed("1111011101011011"),
    signed("0010100000100101"),
    signed("0010000111000000"),
    signed("1111011101100010"),
    signed("0010000111101110"),
    signed("1111111100111000"),
    signed("1111011101100010"),
    signed("0000001111110111"),
    signed("0000101000101110"),
    signed("1101101011011101"),
    signed("1100110011010000"),
    signed("0011001001010010"),
    signed("0010100000100101"),
    signed("1111100110011100"),
    signed("1100011101100001"),
    signed("0000001100000001"),
    signed("0010011001111111"),
    signed("0001000101000010"),
    signed("0000110101111001"),
    signed("0011000011110110"),
    signed("0010010011101111"),
    signed("0000000011001000"),
    signed("1110100111100110"),
    signed("1101000101110111"),
    signed("0010010011101111"),
    signed("0010000111000000"),
    signed("0001001110110000"),
    signed("0001101110001001"));

constant lut_gs2q_data_54 : vector_of_signed16(0 to 63) := 
   (signed("1110100010001111"),
    signed("0010001101011111"),
    signed("0001101100001010"),
    signed("0000001111001111"),
    signed("1100110100100101"),
    signed("1111111100000010"),
    signed("0000001011111110"),
    signed("0000010010100000"),
    signed("0010011010111100"),
    signed("0001110101010110"),
    signed("1110101101000101"),
    signed("1111100110011000"),
    signed("0001111111011000"),
    signed("0010100010001110"),
    signed("0001000100111110"),
    signed("1101100011000110"),
    signed("0000000110001110"),
    signed("1110110010111100"),
    signed("0000001010010011"),
    signed("1111111100000010"),
    signed("0010011100111010"),
    signed("0000110111100001"),
    signed("1100111101111000"),
    signed("0000001110010111"),
    signed("1101101011001111"),
    signed("0001100111001011"),
    signed("0011001111011011"),
    signed("1100110101011010"),
    signed("1101000011101000"),
    signed("1111001111111011"),
    signed("1101001111101011"),
    signed("1110011010001100"),
    signed("1111000000110110"),
    signed("0001100001101100"),
    signed("1110100101111010"),
    signed("0001101001111000"),
    signed("1110100111111100"),
    signed("0010011011000011"),
    signed("0001111111101001"),
    signed("0000010100000111"),
    signed("0010000001101101"),
    signed("1110111011000110"),
    signed("0000010100000111"),
    signed("0000111111011101"),
    signed("1111111110000100"),
    signed("1101100000011001"),
    signed("1100111010010101"),
    signed("0010111110011001"),
    signed("0010101111100100"),
    signed("0000010100101011"),
    signed("1100101000011011"),
    signed("1111010110001111"),
    signed("0010100111111110"),
    signed("0000010011111000"),
    signed("0001011010001101"),
    signed("0011000010001000"),
    signed("0010100001111001"),
    signed("1111010100011000"),
    signed("1110101001001111"),
    signed("1101010000101010"),
    signed("0010100001111001"),
    signed("0001111111101001"),
    signed("0000011000110100"),
    signed("0001100101000000"));

constant lut_gs2q_data_55 : vector_of_signed16(0 to 63) := 
   (signed("1110000011101001"),
    signed("0010010001100100"),
    signed("0001110101100111"),
    signed("0000111000010111"),
    signed("1101000011011001"),
    signed("1111010011001001"),
    signed("1111011000110011"),
    signed("0000110000001101"),
    signed("0010000111010011"),
    signed("0010010110101001"),
    signed("1110010100111111"),
    signed("0000011010011010"),
    signed("0001110010111101"),
    signed("0010100110101110"),
    signed("0001101011100101"),
    signed("1101110010011111"),
    signed("1111010001001100"),
    signed("1110000011011011"),
    signed("0000111000010111"),
    signed("1111010011001001"),
    signed("0010001101100001"),
    signed("0001010010011011"),
    signed("1101001000110101"),
    signed("0001000001110101"),
    signed("1101110010011100"),
    signed("0010000000001000"),
    signed("0011000000110010"),
    signed("1101001010111111"),
    signed("1101010000011011"),
    signed("1110100101010110"),
    signed("1101011110000101"),
    signed("1110010111111101"),
    signed("1110001010111110"),
    signed("0010000111011111"),
    signed("1101111111110100"),
    signed("0001110001100000"),
    signed("1101111101111011"),
    signed("0010010001100011"),
    signed("0001111000111101"),
    signed("0001001001011011"),
    signed("0001111100010111"),
    signed("1110000011010111"),
    signed("0001001001011011"),
    signed("0001100111101011"),
    signed("1111010001010000"),
    signed("1101011011010010"),
    signed("1101001010111111"),
    signed("0010101011100111"),
    signed("0010110101101000"),
    signed("0001000010000100"),
    signed("1100111111010010"),
    signed("1110100101100101"),
    signed("0010101110010101"),
    signed("1111011110000000"),
    signed("0001110100011011"),
    signed("0010110111001011"),
    signed("0010101000110101"),
    signed("1110101001101000"),
    signed("1110100101000000"),
    signed("1101100001011100"),
    signed("0010101000110101"),
    signed("0001111000111101"),
    signed("1111011110000000"),
    signed("0001100000011100"));

constant lut_gs2q_data_56 : vector_of_signed16(0 to 63) := 
   (signed("1101110011101000"),
    signed("0010010010001000"),
    signed("0001111111001110"),
    signed("0001011110110110"),
    signed("1101011011100111"),
    signed("1110101001111110"),
    signed("1110100110010000"),
    signed("0001001111010101"),
    signed("0001110110100000"),
    signed("0010100100101110"),
    signed("1110000110110001"),
    signed("0001001111101110"),
    signed("0001101011101110"),
    signed("0010100001011110"),
    signed("0010000100110100"),
    signed("1110000001101001"),
    signed("1110011110001000"),
    signed("1101100101100001"),
    signed("0001100011000011"),
    signed("1110101001111110"),
    signed("0001111110010111"),
    signed("0001101001000101"),
    signed("1101011100110101"),
    signed("0001101111100100"),
    signed("1101111010010001"),
    signed("0010001010101010"),
    signed("0010100111100000"),
    signed("1101100111111100"),
    signed("1101100100111110"),
    signed("1110000101001001"),
    signed("1101101111011111"),
    signed("1110010001011100"),
    signed("1101100110010010"),
    signed("0010011011110101"),
    signed("1101101001110010"),
    signed("0001111011000110"),
    signed("1101100101010100"),
    signed("0010000100011111"),
    signed("0001110100010101"),
    signed("0001110111101100"),
    signed("0001111001010001"),
    signed("1101011110001001"),
    signed("0001110111101100"),
    signed("0010000100001000"),
    signed("1110100101100000"),
    signed("1101011110111100"),
    signed("1101100011101111"),
    signed("0010010010111011"),
    signed("0010101111001101"),
    signed("0001101010101101"),
    signed("1101011111110111"),
    signed("1110000000010010"),
    signed("0010101001100110"),
    signed("1110101000001001"),
    signed("0010000010100101"),
    signed("0010100011001011"),
    signed("0010100101001100"),
    signed("1110000110011010"),
    signed("1110011010110011"),
    signed("1101110110011100"),
    signed("0010100101001100"),
    signed("0001110100010101"),
    signed("1110100011111101"),
    signed("0001100010001111"));

constant lut_gs2q_data_57 : vector_of_signed16(0 to 63) := 
   (signed("1101110001101100"),
    signed("0010010000110110"),
    signed("0010000101100000"),
    signed("0010000010010010"),
    signed("1101111001100100"),
    signed("1110000000100100"),
    signed("1101110110010101"),
    signed("0001101101000101"),
    signed("0001101001010011"),
    signed("0010011111110101"),
    signed("1110000101011101"),
    signed("0010000100010111"),
    signed("0001101101101001"),
    signed("0010001110100111"),
    signed("0010001111101111"),
    signed("1110001011110000"),
    signed("1101110011101011"),
    signed("1101011011010000"),
    signed("0010000100111100"),
    signed("1110000000100100"),
    signed("0001101111111010"),
    signed("0001111001000001"),
    signed("1101111011010000"),
    signed("0010010001010001"),
    signed("1101111111011011"),
    signed("0010001000001010"),
    signed("0010000111000001"),
    signed("1110000111100100"),
    signed("1110000010010000"),
    signed("1101110101001100"),
    signed("1110000011110010"),
    signed("1110000100110000"),
    signed("1101011010010010"),
    signed("0010011001110011"),
    signed("1101101000110111"),
    signed("0010000111100101"),
    signed("1101011111100110"),
    signed("0001110010000001"),
    signed("0001110100110101"),
    signed("0010011100100111"),
    signed("0001110111010011"),
    signed("1101010011010010"),
    signed("0010011100100111"),
    signed("0010010011111010"),
    signed("1101111011101001"),
    signed("1101101111010100"),
    signed("1110000000100100"),
    signed("0001111000011100"),
    signed("0010011000010001"),
    signed("0010001101101001"),
    signed("1110000101010011"),
    signed("1101101101001110"),
    signed("0010010101100111"),
    signed("1101110100101000"),
    signed("0010000101111001"),
    signed("0010001001000110"),
    signed("0010010010111101"),
    signed("1101101010111110"),
    signed("1110001001000110"),
    signed("1110010000010001"),
    signed("0010010010111101"),
    signed("0001110000011111"),
    signed("1101101101101000"),
    signed("0001101101010000"));

constant lut_gs2q_data_58 : vector_of_signed16(0 to 63) := 
   (signed("1110000010010110"),
    signed("0010000111010110"),
    signed("0010001010001101"),
    signed("0010011110000010"),
    signed("1110100001110110"),
    signed("1101011111110011"),
    signed("1101001111001001"),
    signed("0010001110101110"),
    signed("0001100111110010"),
    signed("0010000010000001"),
    signed("1110001010101101"),
    signed("0010101101111001"),
    signed("0001110110010011"),
    signed("0001110100101110"),
    signed("0010001000100011"),
    signed("1110010101101000"),
    signed("1101001110101011"),
    signed("1101101100010111"),
    signed("0010100010011011"),
    signed("1101011111110011"),
    signed("0001100110101001"),
    signed("0010001000101011"),
    signed("1110011111111101"),
    signed("0010101011000001"),
    signed("1110000011101100"),
    signed("0001110010101110"),
    signed("0001011110101101"),
    signed("1110101110001011"),
    signed("1110100100001001"),
    signed("1101110100111001"),
    signed("1110010010001100"),
    signed("1101111001100001"),
    signed("1101100010010110"),
    signed("0010000111110110"),
    signed("1101110110111011"),
    signed("0010001111000101"),
    signed("1101110000010011"),
    signed("0001100000111101"),
    signed("0001111000000100"),
    signed("0010110010111100"),
    signed("0001111001011110"),
    signed("1101011110001001"),
    signed("0010110010111100"),
    signed("0010001110111010"),
    signed("1101011100111001"),
    signed("1110001010001000"),
    signed("1110100110000010"),
    signed("0001011011001100"),
    signed("0001110111101100"),
    signed("0010100010001110"),
    signed("1110110011010000"),
    signed("1101101000010111"),
    signed("0001111000111011"),
    signed("1101001101111011"),
    signed("0001110111110011"),
    signed("0001100011110010"),
    signed("0001110100101110"),
    signed("1101011110111100"),
    signed("1101111000000101"),
    signed("1110100111000111"),
    signed("0001110100101110"),
    signed("0001110100010101"),
    signed("1101000101110011"),
    signed("0001111010001011"));

constant lut_gs2q_data_59 : vector_of_signed16(0 to 63) := 
   (signed("1110100001101100"),
    signed("0001111101001110"),
    signed("0010001111011110"),
    signed("0010101110010001"),
    signed("1111001011100011"),
    signed("1101000011011001"),
    signed("1100110101110100"),
    signed("0010101011100111"),
    signed("0001101011010111"),
    signed("0001010101001110"),
    signed("1110011100100110"),
    signed("0011001111101000"),
    signed("0010000001110100"),
    signed("0001001110111000"),
    signed("0001101101101011"),
    signed("1110010111111101"),
    signed("1100110111111011"),
    signed("1110010000001011"),
    signed("0010110011110001"),
    signed("1101000011011001"),
    signed("0001100101111100"),
    signed("0010010001100011"),
    signed("1111000110010101"),
    signed("0010110101101000"),
    signed("1110001001000011"),
    signed("0001010011000100"),
    signed("0000101110110000"),
    signed("1111010011001001"),
    signed("1111000110010101"),
    signed("1110000001111110"),
    signed("1110011111100000"),
    signed("1101101010111001"),
    signed("1110000011010111"),
    signed("0001100010000001"),
    signed("1110011000100010"),
    signed("0010010110111110"),
    signed("1110010111110001"),
    signed("0001001010110100"),
    signed("0001111011000100"),
    signed("0010110111101111"),
    signed("0010000001110111"),
    signed("1110000011010111"),
    signed("0010110111101111"),
    signed("0001111100000001"),
    signed("1101000100101110"),
    signed("1110101011101110"),
    signed("1111001011100011"),
    signed("0000111001111010"),
    signed("0001001001011011"),
    signed("0010101110010001"),
    signed("1111100000001010"),
    signed("1101111000100001"),
    signed("0001001110111000"),
    signed("1100110000011000"),
    signed("0001100000000100"),
    signed("0000111011110001"),
    signed("0001001110111000"),
    signed("1101011011010010"),
    signed("1101100011100101"),
    signed("1111000000111001"),
    signed("0001001110111000"),
    signed("0001111000111101"),
    signed("1100101000110001"),
    signed("0010001101100001"));

constant lut_gs2q_data_60 : vector_of_signed16(0 to 63) := 
   (signed("1111001100001000"),
    signed("0001110001111010"),
    signed("0010010010101111"),
    signed("0010110101000011"),
    signed("1111110110010010"),
    signed("1100101111101001"),
    signed("1100101001010011"),
    signed("0011000011010101"),
    signed("0001110100101100"),
    signed("0000011100111011"),
    signed("1110110111110001"),
    signed("0011100100111011"),
    signed("0010001111111100"),
    signed("0000100010010101"),
    signed("0001000100101010"),
    signed("1110010101010000"),
    signed("1100101101111011"),
    signed("1111000011110100"),
    signed("0010111011001000"),
    signed("1100101111101001"),
    signed("0001101011000100"),
    signed("0010010110000111"),
    signed("1111101110011000"),
    signed("0010110100011111"),
    signed("1110001100110110"),
    signed("0000101010010101"),
    signed("1111111101000000"),
    signed("1111110111000111"),
    signed("1111101001011100"),
    signed("1110011101011100"),
    signed("1110101000000110"),
    signed("1101011101010110"),
    signed("1110110110001010"),
    signed("0000101111100001"),
    signed("1111000111001100"),
    signed("0010011100000010"),
    signed("1111001110100000"),
    signed("0000110001110001"),
    signed("0001111111010100"),
    signed("0010101111001111"),
    signed("0010001100101110"),
    signed("1110111011000110"),
    signed("0010101111001111"),
    signed("0001011011000001"),
    signed("1100110110101001"),
    signed("1111010100000011"),
    signed("1111110001010110"),
    signed("0000010111111100"),
    signed("0000010100000111"),
    signed("0010110000001000"),
    signed("0000001011011010"),
    signed("1110011001011000"),
    signed("0000011101011010"),
    signed("1100100000000001"),
    signed("0000111110101000"),
    signed("0000010001010100"),
    signed("0000100010010101"),
    signed("1101100000011001"),
    signed("1101010000110100"),
    signed("1111011011001110"),
    signed("0000100010010101"),
    signed("0001111111101001"),
    signed("1100011010010000"),
    signed("0010100001110110"));

constant lut_gs2q_data_61 : vector_of_signed16(0 to 63) := 
   (signed("1111111100101101"),
    signed("0001100111100100"),
    signed("0010010011110110"),
    signed("0010110011001100"),
    signed("0000011111011101"),
    signed("1100100110011011"),
    signed("1100101001100011"),
    signed("0011010011000000"),
    signed("0010000001001000"),
    signed("1111100000100011"),
    signed("1111011010011010"),
    signed("0011101100001100"),
    signed("0010011101011101"),
    signed("1111110011010001"),
    signed("0000010010100111"),
    signed("1110001110101111"),
    signed("1100110000001000"),
    signed("0000000000000000"),
    signed("0010111001011100"),
    signed("1100100110011011"),
    signed("0001110100011001"),
    signed("0010010110110111"),
    signed("0000010101101111"),
    signed("0010101010010010"),
    signed("1110001110101111"),
    signed("1111111100111000"),
    signed("1111001101100101"),
    signed("0000011000110111"),
    signed("0000001100000001"),
    signed("1111000100101011"),
    signed("1110101011000011"),
    signed("1101010011011010"),
    signed("1111110011001010"),
    signed("1111110111000111"),
    signed("1111111100111000"),
    signed("0010011101011101"),
    signed("0000001100110110"),
    signed("0000010101101111"),
    signed("0010000011111000"),
    signed("0010011101011101"),
    signed("0010010111101011"),
    signed("1111111100111000"),
    signed("0010011101011101"),
    signed("0000101111010011"),
    signed("1100110011010000"),
    signed("0000000000000000"),
    signed("0000010101101111"),
    signed("1111110110010010"),
    signed("1111011101100010"),
    signed("0010101001011110"),
    signed("0000110010011011"),
    signed("1111000110111111"),
    signed("1111101001100100"),
    signed("1100011101100001"),
    signed("0000010110011100"),
    signed("1111100111001001"),
    signed("1111110011010001"),
    signed("1101101011011101"),
    signed("1101000011000111"),
    signed("1111110110010010"),
    signed("1111110011010001"),
    signed("0010000111000000"),
    signed("1100011010011001"),
    signed("0010110011001100"));

constant lut_gs2q_data_62 : vector_of_signed16(0 to 63) := 
   (signed("0000101101110010"),
    signed("0001100000011000"),
    signed("0010010010101111"),
    signed("0010101010010000"),
    signed("0001000100100011"),
    signed("1100101000111111"),
    signed("1100110101011010"),
    signed("0011010111110110"),
    signed("0010001101010101"),
    signed("1110101000010000"),
    signed("0000000010010000"),
    signed("0011100100111011"),
    signed("0010100110110101"),
    signed("1111000110010011"),
    signed("1111011101110101"),
    signed("1110000110001011"),
    signed("1100111100111111"),
    signed("0000111100001100"),
    signed("0010110000010101"),
    signed("1100101000111111"),
    signed("0001111111100101"),
    signed("0010010100011100"),
    signed("0000111010001011"),
    signed("0010011010101000"),
    signed("1110001110100110"),
    signed("1111001111100110"),
    signed("1110100100101010"),
    signed("0000110111100001"),
    signed("0000101100110101"),
    signed("1111110100000010"),
    signed("1110101000000110"),
    signed("1101001111100100"),
    signed("0000110001100000"),
    signed("1111000000010010"),
    signed("0000110010101111"),
    signed("0010011010101111"),
    signed("0001001001110110"),
    signed("1111110110110010"),
    signed("0010000111101111"),
    signed("0010000111100001"),
    signed("0010011111111011"),
    signed("0000111110110110"),
    signed("0010000111100001"),
    signed("1111111101001111"),
    signed("1100111010010101"),
    signed("0000101011111101"),
    signed("0000110111001101"),
    signed("1111010101110010"),
    signed("1110101011111111"),
    signed("0010011100111010"),
    signed("0001010010111011"),
    signed("1111111100000101"),
    signed("1110111000111101"),
    signed("1100101000011011"),
    signed("1111101011000001"),
    signed("1111000000000101"),
    signed("1111000110010011"),
    signed("1101111001000011"),
    signed("1100111101100111"),
    signed("0000010010100000"),
    signed("1111000110010011"),
    signed("0010001101011111"),
    signed("1100101000000111"),
    signed("0010111101011110"));

constant lut_gs2q_data_63 : vector_of_signed16(0 to 63) := 
   (signed("0001011001100111"),
    signed("0001011110010110"),
    signed("0010001111011110"),
    signed("0010011100011011"),
    signed("0001100011011011"),
    signed("1100110111111011"),
    signed("1101001010111111"),
    signed("0011001111101100"),
    signed("0010010101110100"),
    signed("1101111011110101"),
    signed("0000101100101010"),
    signed("0011001111101000"),
    signed("0010101000110101"),
    signed("1110011111111100"),
    signed("1110101100111001"),
    signed("1101111101100101"),
    signed("1101010010010011"),
    signed("0001101111110101"),
    signed("0010100001111011"),
    signed("1100110111111011"),
    signed("0010001010000001"),
    signed("0010001111101011"),
    signed("0001011001101110"),
    signed("0010001001011010"),
    signed("1110001100011111"),
    signed("1110100111011100"),
    signed("1110000110000101"),
    signed("0001010010011011"),
    signed("0001001010110100"),
    signed("0000100111001101"),
    signed("1110011111100000"),
    signed("1101010011110101"),
    signed("0001101000001111"),
    signed("1110010010010101"),
    signed("0001100001111110"),
    signed("0010010011101010"),
    signed("0001111100101001"),
    signed("1111010101001111"),
    signed("0010001001111110"),
    signed("0001110010111010"),
    signed("0010100010100111"),
    signed("0001110111001001"),
    signed("0001110010111010"),
    signed("1111001001101001"),
    signed("1101001010111111"),
    signed("0001010100010010"),
    signed("0001010100100001"),
    signed("1110110111001100"),
    signed("1110000101010100"),
    signed("0010001101100001"),
    signed("0001101011000001"),
    signed("0000110010111011"),
    signed("1110010001000010"),
    signed("1100111111010010"),
    signed("1111000000000011"),
    signed("1110011110101011"),
    signed("1110011111111100"),
    signed("1110000101101111"),
    signed("1101000010110101"),
    signed("0000110000001101"),
    signed("1110011111111100"),
    signed("0010010001100100"),
    signed("1101000001011000"),
    signed("0010111101001011"));

constant lut_gs2q_data_64 : vector_of_signed16(0 to 63) := 
   (signed("0001111011000110"),
    signed("0001100010101101"),
    signed("0010001010001101"),
    signed("0010001100000111"),
    signed("0001111010100100"),
    signed("1101010010111000"),
    signed("1101100111111100"),
    signed("0010111001011101"),
    signed("0010010111100000"),
    signed("1101100001100101"),
    signed("0001010110110010"),
    signed("0010101101111001"),
    signed("0010100001000000"),
    signed("1110000100000000"),
    signed("1110000101111010"),
    signed("1101110110110000"),
    signed("1101101101100011"),
    signed("0010010011101001"),
    signed("0010010000100001"),
    signed("1101010010111000"),
    signed("0010010001011000"),
    signed("0010001001011101"),
    signed("0001110010111010"),
    signed("0001111010001111"),
    signed("1110001000101101"),
    signed("1110001000111000"),
    signed("1101110100110100"),
    signed("0001101001000101"),
    signed("0001100101001010"),
    signed("0001011001110000"),
    signed("1110010010001100"),
    signed("1101100001100000"),
    signed("0010001111101101"),
    signed("1101110011010001"),
    signed("0010000100101011"),
    signed("0010001000001101"),
    signed("0010011101101010"),
    signed("1110110001111001"),
    signed("0010001010000000"),
    signed("0001100100010110"),
    signed("0010011101010101"),
    signed("0010011101011101"),
    signed("0001100100010110"),
    signed("1110011001001011"),
    signed("1101100011101111"),
    signed("0001110101111000"),
    signed("0001101100110100"),
    signed("1110011011010000"),
    signed("1101101110001100"),
    signed("0001111110010111"),
    signed("0001111001001111"),
    signed("0001100110000001"),
    signed("1101110110010000"),
    signed("1101011111110111"),
    signed("1110011001000010"),
    signed("1110000100111110"),
    signed("1110000100000000"),
    signed("1110001110101010"),
    signed("1101010100001110"),
    signed("0001001111010101"),
    signed("1110000100000000"),
    signed("0010010010001000"),
    signed("1101100011100110"),
    signed("0010101111111110"));

